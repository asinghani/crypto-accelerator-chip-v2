magic
tech sky130A
magscale 1 2
timestamp 1636415114
<< obsli1 >>
rect 1104 1309 310868 311729
<< obsm1 >>
rect 1104 1303 311130 311760
<< metal2 >>
rect 1306 313367 1362 314167
rect 3974 313367 4030 314167
rect 6734 313367 6790 314167
rect 9494 313367 9550 314167
rect 12254 313367 12310 314167
rect 14922 313367 14978 314167
rect 17682 313367 17738 314167
rect 20442 313367 20498 314167
rect 23202 313367 23258 314167
rect 25870 313367 25926 314167
rect 28630 313367 28686 314167
rect 31390 313367 31446 314167
rect 34150 313367 34206 314167
rect 36818 313367 36874 314167
rect 39578 313367 39634 314167
rect 42338 313367 42394 314167
rect 45098 313367 45154 314167
rect 47766 313367 47822 314167
rect 50526 313367 50582 314167
rect 53286 313367 53342 314167
rect 56046 313367 56102 314167
rect 58714 313367 58770 314167
rect 61474 313367 61530 314167
rect 64234 313367 64290 314167
rect 66994 313367 67050 314167
rect 69662 313367 69718 314167
rect 72422 313367 72478 314167
rect 75182 313367 75238 314167
rect 77942 313367 77998 314167
rect 80610 313367 80666 314167
rect 83370 313367 83426 314167
rect 86130 313367 86186 314167
rect 88890 313367 88946 314167
rect 91558 313367 91614 314167
rect 94318 313367 94374 314167
rect 97078 313367 97134 314167
rect 99838 313367 99894 314167
rect 102506 313367 102562 314167
rect 105266 313367 105322 314167
rect 108026 313367 108082 314167
rect 110786 313367 110842 314167
rect 113454 313367 113510 314167
rect 116214 313367 116270 314167
rect 118974 313367 119030 314167
rect 121734 313367 121790 314167
rect 124402 313367 124458 314167
rect 127162 313367 127218 314167
rect 129922 313367 129978 314167
rect 132682 313367 132738 314167
rect 135350 313367 135406 314167
rect 138110 313367 138166 314167
rect 140870 313367 140926 314167
rect 143630 313367 143686 314167
rect 146298 313367 146354 314167
rect 149058 313367 149114 314167
rect 151818 313367 151874 314167
rect 154578 313367 154634 314167
rect 157338 313367 157394 314167
rect 160006 313367 160062 314167
rect 162766 313367 162822 314167
rect 165526 313367 165582 314167
rect 168286 313367 168342 314167
rect 170954 313367 171010 314167
rect 173714 313367 173770 314167
rect 176474 313367 176530 314167
rect 179234 313367 179290 314167
rect 181902 313367 181958 314167
rect 184662 313367 184718 314167
rect 187422 313367 187478 314167
rect 190182 313367 190238 314167
rect 192850 313367 192906 314167
rect 195610 313367 195666 314167
rect 198370 313367 198426 314167
rect 201130 313367 201186 314167
rect 203798 313367 203854 314167
rect 206558 313367 206614 314167
rect 209318 313367 209374 314167
rect 212078 313367 212134 314167
rect 214746 313367 214802 314167
rect 217506 313367 217562 314167
rect 220266 313367 220322 314167
rect 223026 313367 223082 314167
rect 225694 313367 225750 314167
rect 228454 313367 228510 314167
rect 231214 313367 231270 314167
rect 233974 313367 234030 314167
rect 236642 313367 236698 314167
rect 239402 313367 239458 314167
rect 242162 313367 242218 314167
rect 244922 313367 244978 314167
rect 247590 313367 247646 314167
rect 250350 313367 250406 314167
rect 253110 313367 253166 314167
rect 255870 313367 255926 314167
rect 258538 313367 258594 314167
rect 261298 313367 261354 314167
rect 264058 313367 264114 314167
rect 266818 313367 266874 314167
rect 269486 313367 269542 314167
rect 272246 313367 272302 314167
rect 275006 313367 275062 314167
rect 277766 313367 277822 314167
rect 280434 313367 280490 314167
rect 283194 313367 283250 314167
rect 285954 313367 286010 314167
rect 288714 313367 288770 314167
rect 291382 313367 291438 314167
rect 294142 313367 294198 314167
rect 296902 313367 296958 314167
rect 299662 313367 299718 314167
rect 302330 313367 302386 314167
rect 305090 313367 305146 314167
rect 307850 313367 307906 314167
rect 310610 313367 310666 314167
rect 294 0 350 800
rect 846 0 902 800
rect 1490 0 1546 800
rect 2134 0 2190 800
rect 2778 0 2834 800
rect 3422 0 3478 800
rect 4066 0 4122 800
rect 4710 0 4766 800
rect 5354 0 5410 800
rect 5998 0 6054 800
rect 6642 0 6698 800
rect 7286 0 7342 800
rect 7930 0 7986 800
rect 8482 0 8538 800
rect 9126 0 9182 800
rect 9770 0 9826 800
rect 10414 0 10470 800
rect 11058 0 11114 800
rect 11702 0 11758 800
rect 12346 0 12402 800
rect 12990 0 13046 800
rect 13634 0 13690 800
rect 14278 0 14334 800
rect 14922 0 14978 800
rect 15566 0 15622 800
rect 16210 0 16266 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25042 0 25098 800
rect 25686 0 25742 800
rect 26330 0 26386 800
rect 26974 0 27030 800
rect 27618 0 27674 800
rect 28262 0 28318 800
rect 28906 0 28962 800
rect 29550 0 29606 800
rect 30194 0 30250 800
rect 30838 0 30894 800
rect 31482 0 31538 800
rect 32126 0 32182 800
rect 32770 0 32826 800
rect 33322 0 33378 800
rect 33966 0 34022 800
rect 34610 0 34666 800
rect 35254 0 35310 800
rect 35898 0 35954 800
rect 36542 0 36598 800
rect 37186 0 37242 800
rect 37830 0 37886 800
rect 38474 0 38530 800
rect 39118 0 39174 800
rect 39762 0 39818 800
rect 40406 0 40462 800
rect 41050 0 41106 800
rect 41602 0 41658 800
rect 42246 0 42302 800
rect 42890 0 42946 800
rect 43534 0 43590 800
rect 44178 0 44234 800
rect 44822 0 44878 800
rect 45466 0 45522 800
rect 46110 0 46166 800
rect 46754 0 46810 800
rect 47398 0 47454 800
rect 48042 0 48098 800
rect 48686 0 48742 800
rect 49330 0 49386 800
rect 49882 0 49938 800
rect 50526 0 50582 800
rect 51170 0 51226 800
rect 51814 0 51870 800
rect 52458 0 52514 800
rect 53102 0 53158 800
rect 53746 0 53802 800
rect 54390 0 54446 800
rect 55034 0 55090 800
rect 55678 0 55734 800
rect 56322 0 56378 800
rect 56966 0 57022 800
rect 57610 0 57666 800
rect 58162 0 58218 800
rect 58806 0 58862 800
rect 59450 0 59506 800
rect 60094 0 60150 800
rect 60738 0 60794 800
rect 61382 0 61438 800
rect 62026 0 62082 800
rect 62670 0 62726 800
rect 63314 0 63370 800
rect 63958 0 64014 800
rect 64602 0 64658 800
rect 65246 0 65302 800
rect 65890 0 65946 800
rect 66442 0 66498 800
rect 67086 0 67142 800
rect 67730 0 67786 800
rect 68374 0 68430 800
rect 69018 0 69074 800
rect 69662 0 69718 800
rect 70306 0 70362 800
rect 70950 0 71006 800
rect 71594 0 71650 800
rect 72238 0 72294 800
rect 72882 0 72938 800
rect 73526 0 73582 800
rect 74170 0 74226 800
rect 74722 0 74778 800
rect 75366 0 75422 800
rect 76010 0 76066 800
rect 76654 0 76710 800
rect 77298 0 77354 800
rect 77942 0 77998 800
rect 78586 0 78642 800
rect 79230 0 79286 800
rect 79874 0 79930 800
rect 80518 0 80574 800
rect 81162 0 81218 800
rect 81806 0 81862 800
rect 82358 0 82414 800
rect 83002 0 83058 800
rect 83646 0 83702 800
rect 84290 0 84346 800
rect 84934 0 84990 800
rect 85578 0 85634 800
rect 86222 0 86278 800
rect 86866 0 86922 800
rect 87510 0 87566 800
rect 88154 0 88210 800
rect 88798 0 88854 800
rect 89442 0 89498 800
rect 90086 0 90142 800
rect 90638 0 90694 800
rect 91282 0 91338 800
rect 91926 0 91982 800
rect 92570 0 92626 800
rect 93214 0 93270 800
rect 93858 0 93914 800
rect 94502 0 94558 800
rect 95146 0 95202 800
rect 95790 0 95846 800
rect 96434 0 96490 800
rect 97078 0 97134 800
rect 97722 0 97778 800
rect 98366 0 98422 800
rect 98918 0 98974 800
rect 99562 0 99618 800
rect 100206 0 100262 800
rect 100850 0 100906 800
rect 101494 0 101550 800
rect 102138 0 102194 800
rect 102782 0 102838 800
rect 103426 0 103482 800
rect 104070 0 104126 800
rect 104714 0 104770 800
rect 105358 0 105414 800
rect 106002 0 106058 800
rect 106646 0 106702 800
rect 107198 0 107254 800
rect 107842 0 107898 800
rect 108486 0 108542 800
rect 109130 0 109186 800
rect 109774 0 109830 800
rect 110418 0 110474 800
rect 111062 0 111118 800
rect 111706 0 111762 800
rect 112350 0 112406 800
rect 112994 0 113050 800
rect 113638 0 113694 800
rect 114282 0 114338 800
rect 114926 0 114982 800
rect 115478 0 115534 800
rect 116122 0 116178 800
rect 116766 0 116822 800
rect 117410 0 117466 800
rect 118054 0 118110 800
rect 118698 0 118754 800
rect 119342 0 119398 800
rect 119986 0 120042 800
rect 120630 0 120686 800
rect 121274 0 121330 800
rect 121918 0 121974 800
rect 122562 0 122618 800
rect 123206 0 123262 800
rect 123758 0 123814 800
rect 124402 0 124458 800
rect 125046 0 125102 800
rect 125690 0 125746 800
rect 126334 0 126390 800
rect 126978 0 127034 800
rect 127622 0 127678 800
rect 128266 0 128322 800
rect 128910 0 128966 800
rect 129554 0 129610 800
rect 130198 0 130254 800
rect 130842 0 130898 800
rect 131486 0 131542 800
rect 132038 0 132094 800
rect 132682 0 132738 800
rect 133326 0 133382 800
rect 133970 0 134026 800
rect 134614 0 134670 800
rect 135258 0 135314 800
rect 135902 0 135958 800
rect 136546 0 136602 800
rect 137190 0 137246 800
rect 137834 0 137890 800
rect 138478 0 138534 800
rect 139122 0 139178 800
rect 139766 0 139822 800
rect 140318 0 140374 800
rect 140962 0 141018 800
rect 141606 0 141662 800
rect 142250 0 142306 800
rect 142894 0 142950 800
rect 143538 0 143594 800
rect 144182 0 144238 800
rect 144826 0 144882 800
rect 145470 0 145526 800
rect 146114 0 146170 800
rect 146758 0 146814 800
rect 147402 0 147458 800
rect 148046 0 148102 800
rect 148598 0 148654 800
rect 149242 0 149298 800
rect 149886 0 149942 800
rect 150530 0 150586 800
rect 151174 0 151230 800
rect 151818 0 151874 800
rect 152462 0 152518 800
rect 153106 0 153162 800
rect 153750 0 153806 800
rect 154394 0 154450 800
rect 155038 0 155094 800
rect 155682 0 155738 800
rect 156326 0 156382 800
rect 156878 0 156934 800
rect 157522 0 157578 800
rect 158166 0 158222 800
rect 158810 0 158866 800
rect 159454 0 159510 800
rect 160098 0 160154 800
rect 160742 0 160798 800
rect 161386 0 161442 800
rect 162030 0 162086 800
rect 162674 0 162730 800
rect 163318 0 163374 800
rect 163962 0 164018 800
rect 164514 0 164570 800
rect 165158 0 165214 800
rect 165802 0 165858 800
rect 166446 0 166502 800
rect 167090 0 167146 800
rect 167734 0 167790 800
rect 168378 0 168434 800
rect 169022 0 169078 800
rect 169666 0 169722 800
rect 170310 0 170366 800
rect 170954 0 171010 800
rect 171598 0 171654 800
rect 172242 0 172298 800
rect 172794 0 172850 800
rect 173438 0 173494 800
rect 174082 0 174138 800
rect 174726 0 174782 800
rect 175370 0 175426 800
rect 176014 0 176070 800
rect 176658 0 176714 800
rect 177302 0 177358 800
rect 177946 0 178002 800
rect 178590 0 178646 800
rect 179234 0 179290 800
rect 179878 0 179934 800
rect 180522 0 180578 800
rect 181074 0 181130 800
rect 181718 0 181774 800
rect 182362 0 182418 800
rect 183006 0 183062 800
rect 183650 0 183706 800
rect 184294 0 184350 800
rect 184938 0 184994 800
rect 185582 0 185638 800
rect 186226 0 186282 800
rect 186870 0 186926 800
rect 187514 0 187570 800
rect 188158 0 188214 800
rect 188802 0 188858 800
rect 189354 0 189410 800
rect 189998 0 190054 800
rect 190642 0 190698 800
rect 191286 0 191342 800
rect 191930 0 191986 800
rect 192574 0 192630 800
rect 193218 0 193274 800
rect 193862 0 193918 800
rect 194506 0 194562 800
rect 195150 0 195206 800
rect 195794 0 195850 800
rect 196438 0 196494 800
rect 197082 0 197138 800
rect 197634 0 197690 800
rect 198278 0 198334 800
rect 198922 0 198978 800
rect 199566 0 199622 800
rect 200210 0 200266 800
rect 200854 0 200910 800
rect 201498 0 201554 800
rect 202142 0 202198 800
rect 202786 0 202842 800
rect 203430 0 203486 800
rect 204074 0 204130 800
rect 204718 0 204774 800
rect 205362 0 205418 800
rect 205914 0 205970 800
rect 206558 0 206614 800
rect 207202 0 207258 800
rect 207846 0 207902 800
rect 208490 0 208546 800
rect 209134 0 209190 800
rect 209778 0 209834 800
rect 210422 0 210478 800
rect 211066 0 211122 800
rect 211710 0 211766 800
rect 212354 0 212410 800
rect 212998 0 213054 800
rect 213642 0 213698 800
rect 214194 0 214250 800
rect 214838 0 214894 800
rect 215482 0 215538 800
rect 216126 0 216182 800
rect 216770 0 216826 800
rect 217414 0 217470 800
rect 218058 0 218114 800
rect 218702 0 218758 800
rect 219346 0 219402 800
rect 219990 0 220046 800
rect 220634 0 220690 800
rect 221278 0 221334 800
rect 221922 0 221978 800
rect 222474 0 222530 800
rect 223118 0 223174 800
rect 223762 0 223818 800
rect 224406 0 224462 800
rect 225050 0 225106 800
rect 225694 0 225750 800
rect 226338 0 226394 800
rect 226982 0 227038 800
rect 227626 0 227682 800
rect 228270 0 228326 800
rect 228914 0 228970 800
rect 229558 0 229614 800
rect 230202 0 230258 800
rect 230754 0 230810 800
rect 231398 0 231454 800
rect 232042 0 232098 800
rect 232686 0 232742 800
rect 233330 0 233386 800
rect 233974 0 234030 800
rect 234618 0 234674 800
rect 235262 0 235318 800
rect 235906 0 235962 800
rect 236550 0 236606 800
rect 237194 0 237250 800
rect 237838 0 237894 800
rect 238390 0 238446 800
rect 239034 0 239090 800
rect 239678 0 239734 800
rect 240322 0 240378 800
rect 240966 0 241022 800
rect 241610 0 241666 800
rect 242254 0 242310 800
rect 242898 0 242954 800
rect 243542 0 243598 800
rect 244186 0 244242 800
rect 244830 0 244886 800
rect 245474 0 245530 800
rect 246118 0 246174 800
rect 246670 0 246726 800
rect 247314 0 247370 800
rect 247958 0 248014 800
rect 248602 0 248658 800
rect 249246 0 249302 800
rect 249890 0 249946 800
rect 250534 0 250590 800
rect 251178 0 251234 800
rect 251822 0 251878 800
rect 252466 0 252522 800
rect 253110 0 253166 800
rect 253754 0 253810 800
rect 254398 0 254454 800
rect 254950 0 255006 800
rect 255594 0 255650 800
rect 256238 0 256294 800
rect 256882 0 256938 800
rect 257526 0 257582 800
rect 258170 0 258226 800
rect 258814 0 258870 800
rect 259458 0 259514 800
rect 260102 0 260158 800
rect 260746 0 260802 800
rect 261390 0 261446 800
rect 262034 0 262090 800
rect 262678 0 262734 800
rect 263230 0 263286 800
rect 263874 0 263930 800
rect 264518 0 264574 800
rect 265162 0 265218 800
rect 265806 0 265862 800
rect 266450 0 266506 800
rect 267094 0 267150 800
rect 267738 0 267794 800
rect 268382 0 268438 800
rect 269026 0 269082 800
rect 269670 0 269726 800
rect 270314 0 270370 800
rect 270958 0 271014 800
rect 271510 0 271566 800
rect 272154 0 272210 800
rect 272798 0 272854 800
rect 273442 0 273498 800
rect 274086 0 274142 800
rect 274730 0 274786 800
rect 275374 0 275430 800
rect 276018 0 276074 800
rect 276662 0 276718 800
rect 277306 0 277362 800
rect 277950 0 278006 800
rect 278594 0 278650 800
rect 279238 0 279294 800
rect 279790 0 279846 800
rect 280434 0 280490 800
rect 281078 0 281134 800
rect 281722 0 281778 800
rect 282366 0 282422 800
rect 283010 0 283066 800
rect 283654 0 283710 800
rect 284298 0 284354 800
rect 284942 0 284998 800
rect 285586 0 285642 800
rect 286230 0 286286 800
rect 286874 0 286930 800
rect 287518 0 287574 800
rect 288070 0 288126 800
rect 288714 0 288770 800
rect 289358 0 289414 800
rect 290002 0 290058 800
rect 290646 0 290702 800
rect 291290 0 291346 800
rect 291934 0 291990 800
rect 292578 0 292634 800
rect 293222 0 293278 800
rect 293866 0 293922 800
rect 294510 0 294566 800
rect 295154 0 295210 800
rect 295798 0 295854 800
rect 296350 0 296406 800
rect 296994 0 297050 800
rect 297638 0 297694 800
rect 298282 0 298338 800
rect 298926 0 298982 800
rect 299570 0 299626 800
rect 300214 0 300270 800
rect 300858 0 300914 800
rect 301502 0 301558 800
rect 302146 0 302202 800
rect 302790 0 302846 800
rect 303434 0 303490 800
rect 304078 0 304134 800
rect 304630 0 304686 800
rect 305274 0 305330 800
rect 305918 0 305974 800
rect 306562 0 306618 800
rect 307206 0 307262 800
rect 307850 0 307906 800
rect 308494 0 308550 800
rect 309138 0 309194 800
rect 309782 0 309838 800
rect 310426 0 310482 800
rect 311070 0 311126 800
rect 311714 0 311770 800
<< obsm2 >>
rect 294 313311 1250 313426
rect 1418 313311 3918 313426
rect 4086 313311 6678 313426
rect 6846 313311 9438 313426
rect 9606 313311 12198 313426
rect 12366 313311 14866 313426
rect 15034 313311 17626 313426
rect 17794 313311 20386 313426
rect 20554 313311 23146 313426
rect 23314 313311 25814 313426
rect 25982 313311 28574 313426
rect 28742 313311 31334 313426
rect 31502 313311 34094 313426
rect 34262 313311 36762 313426
rect 36930 313311 39522 313426
rect 39690 313311 42282 313426
rect 42450 313311 45042 313426
rect 45210 313311 47710 313426
rect 47878 313311 50470 313426
rect 50638 313311 53230 313426
rect 53398 313311 55990 313426
rect 56158 313311 58658 313426
rect 58826 313311 61418 313426
rect 61586 313311 64178 313426
rect 64346 313311 66938 313426
rect 67106 313311 69606 313426
rect 69774 313311 72366 313426
rect 72534 313311 75126 313426
rect 75294 313311 77886 313426
rect 78054 313311 80554 313426
rect 80722 313311 83314 313426
rect 83482 313311 86074 313426
rect 86242 313311 88834 313426
rect 89002 313311 91502 313426
rect 91670 313311 94262 313426
rect 94430 313311 97022 313426
rect 97190 313311 99782 313426
rect 99950 313311 102450 313426
rect 102618 313311 105210 313426
rect 105378 313311 107970 313426
rect 108138 313311 110730 313426
rect 110898 313311 113398 313426
rect 113566 313311 116158 313426
rect 116326 313311 118918 313426
rect 119086 313311 121678 313426
rect 121846 313311 124346 313426
rect 124514 313311 127106 313426
rect 127274 313311 129866 313426
rect 130034 313311 132626 313426
rect 132794 313311 135294 313426
rect 135462 313311 138054 313426
rect 138222 313311 140814 313426
rect 140982 313311 143574 313426
rect 143742 313311 146242 313426
rect 146410 313311 149002 313426
rect 149170 313311 151762 313426
rect 151930 313311 154522 313426
rect 154690 313311 157282 313426
rect 157450 313311 159950 313426
rect 160118 313311 162710 313426
rect 162878 313311 165470 313426
rect 165638 313311 168230 313426
rect 168398 313311 170898 313426
rect 171066 313311 173658 313426
rect 173826 313311 176418 313426
rect 176586 313311 179178 313426
rect 179346 313311 181846 313426
rect 182014 313311 184606 313426
rect 184774 313311 187366 313426
rect 187534 313311 190126 313426
rect 190294 313311 192794 313426
rect 192962 313311 195554 313426
rect 195722 313311 198314 313426
rect 198482 313311 201074 313426
rect 201242 313311 203742 313426
rect 203910 313311 206502 313426
rect 206670 313311 209262 313426
rect 209430 313311 212022 313426
rect 212190 313311 214690 313426
rect 214858 313311 217450 313426
rect 217618 313311 220210 313426
rect 220378 313311 222970 313426
rect 223138 313311 225638 313426
rect 225806 313311 228398 313426
rect 228566 313311 231158 313426
rect 231326 313311 233918 313426
rect 234086 313311 236586 313426
rect 236754 313311 239346 313426
rect 239514 313311 242106 313426
rect 242274 313311 244866 313426
rect 245034 313311 247534 313426
rect 247702 313311 250294 313426
rect 250462 313311 253054 313426
rect 253222 313311 255814 313426
rect 255982 313311 258482 313426
rect 258650 313311 261242 313426
rect 261410 313311 264002 313426
rect 264170 313311 266762 313426
rect 266930 313311 269430 313426
rect 269598 313311 272190 313426
rect 272358 313311 274950 313426
rect 275118 313311 277710 313426
rect 277878 313311 280378 313426
rect 280546 313311 283138 313426
rect 283306 313311 285898 313426
rect 286066 313311 288658 313426
rect 288826 313311 291326 313426
rect 291494 313311 294086 313426
rect 294254 313311 296846 313426
rect 297014 313311 299606 313426
rect 299774 313311 302274 313426
rect 302442 313311 305034 313426
rect 305202 313311 307794 313426
rect 307962 313311 310554 313426
rect 310722 313311 311124 313426
rect 294 856 311124 313311
rect 406 734 790 856
rect 958 734 1434 856
rect 1602 734 2078 856
rect 2246 734 2722 856
rect 2890 734 3366 856
rect 3534 734 4010 856
rect 4178 734 4654 856
rect 4822 734 5298 856
rect 5466 734 5942 856
rect 6110 734 6586 856
rect 6754 734 7230 856
rect 7398 734 7874 856
rect 8042 734 8426 856
rect 8594 734 9070 856
rect 9238 734 9714 856
rect 9882 734 10358 856
rect 10526 734 11002 856
rect 11170 734 11646 856
rect 11814 734 12290 856
rect 12458 734 12934 856
rect 13102 734 13578 856
rect 13746 734 14222 856
rect 14390 734 14866 856
rect 15034 734 15510 856
rect 15678 734 16154 856
rect 16322 734 16706 856
rect 16874 734 17350 856
rect 17518 734 17994 856
rect 18162 734 18638 856
rect 18806 734 19282 856
rect 19450 734 19926 856
rect 20094 734 20570 856
rect 20738 734 21214 856
rect 21382 734 21858 856
rect 22026 734 22502 856
rect 22670 734 23146 856
rect 23314 734 23790 856
rect 23958 734 24434 856
rect 24602 734 24986 856
rect 25154 734 25630 856
rect 25798 734 26274 856
rect 26442 734 26918 856
rect 27086 734 27562 856
rect 27730 734 28206 856
rect 28374 734 28850 856
rect 29018 734 29494 856
rect 29662 734 30138 856
rect 30306 734 30782 856
rect 30950 734 31426 856
rect 31594 734 32070 856
rect 32238 734 32714 856
rect 32882 734 33266 856
rect 33434 734 33910 856
rect 34078 734 34554 856
rect 34722 734 35198 856
rect 35366 734 35842 856
rect 36010 734 36486 856
rect 36654 734 37130 856
rect 37298 734 37774 856
rect 37942 734 38418 856
rect 38586 734 39062 856
rect 39230 734 39706 856
rect 39874 734 40350 856
rect 40518 734 40994 856
rect 41162 734 41546 856
rect 41714 734 42190 856
rect 42358 734 42834 856
rect 43002 734 43478 856
rect 43646 734 44122 856
rect 44290 734 44766 856
rect 44934 734 45410 856
rect 45578 734 46054 856
rect 46222 734 46698 856
rect 46866 734 47342 856
rect 47510 734 47986 856
rect 48154 734 48630 856
rect 48798 734 49274 856
rect 49442 734 49826 856
rect 49994 734 50470 856
rect 50638 734 51114 856
rect 51282 734 51758 856
rect 51926 734 52402 856
rect 52570 734 53046 856
rect 53214 734 53690 856
rect 53858 734 54334 856
rect 54502 734 54978 856
rect 55146 734 55622 856
rect 55790 734 56266 856
rect 56434 734 56910 856
rect 57078 734 57554 856
rect 57722 734 58106 856
rect 58274 734 58750 856
rect 58918 734 59394 856
rect 59562 734 60038 856
rect 60206 734 60682 856
rect 60850 734 61326 856
rect 61494 734 61970 856
rect 62138 734 62614 856
rect 62782 734 63258 856
rect 63426 734 63902 856
rect 64070 734 64546 856
rect 64714 734 65190 856
rect 65358 734 65834 856
rect 66002 734 66386 856
rect 66554 734 67030 856
rect 67198 734 67674 856
rect 67842 734 68318 856
rect 68486 734 68962 856
rect 69130 734 69606 856
rect 69774 734 70250 856
rect 70418 734 70894 856
rect 71062 734 71538 856
rect 71706 734 72182 856
rect 72350 734 72826 856
rect 72994 734 73470 856
rect 73638 734 74114 856
rect 74282 734 74666 856
rect 74834 734 75310 856
rect 75478 734 75954 856
rect 76122 734 76598 856
rect 76766 734 77242 856
rect 77410 734 77886 856
rect 78054 734 78530 856
rect 78698 734 79174 856
rect 79342 734 79818 856
rect 79986 734 80462 856
rect 80630 734 81106 856
rect 81274 734 81750 856
rect 81918 734 82302 856
rect 82470 734 82946 856
rect 83114 734 83590 856
rect 83758 734 84234 856
rect 84402 734 84878 856
rect 85046 734 85522 856
rect 85690 734 86166 856
rect 86334 734 86810 856
rect 86978 734 87454 856
rect 87622 734 88098 856
rect 88266 734 88742 856
rect 88910 734 89386 856
rect 89554 734 90030 856
rect 90198 734 90582 856
rect 90750 734 91226 856
rect 91394 734 91870 856
rect 92038 734 92514 856
rect 92682 734 93158 856
rect 93326 734 93802 856
rect 93970 734 94446 856
rect 94614 734 95090 856
rect 95258 734 95734 856
rect 95902 734 96378 856
rect 96546 734 97022 856
rect 97190 734 97666 856
rect 97834 734 98310 856
rect 98478 734 98862 856
rect 99030 734 99506 856
rect 99674 734 100150 856
rect 100318 734 100794 856
rect 100962 734 101438 856
rect 101606 734 102082 856
rect 102250 734 102726 856
rect 102894 734 103370 856
rect 103538 734 104014 856
rect 104182 734 104658 856
rect 104826 734 105302 856
rect 105470 734 105946 856
rect 106114 734 106590 856
rect 106758 734 107142 856
rect 107310 734 107786 856
rect 107954 734 108430 856
rect 108598 734 109074 856
rect 109242 734 109718 856
rect 109886 734 110362 856
rect 110530 734 111006 856
rect 111174 734 111650 856
rect 111818 734 112294 856
rect 112462 734 112938 856
rect 113106 734 113582 856
rect 113750 734 114226 856
rect 114394 734 114870 856
rect 115038 734 115422 856
rect 115590 734 116066 856
rect 116234 734 116710 856
rect 116878 734 117354 856
rect 117522 734 117998 856
rect 118166 734 118642 856
rect 118810 734 119286 856
rect 119454 734 119930 856
rect 120098 734 120574 856
rect 120742 734 121218 856
rect 121386 734 121862 856
rect 122030 734 122506 856
rect 122674 734 123150 856
rect 123318 734 123702 856
rect 123870 734 124346 856
rect 124514 734 124990 856
rect 125158 734 125634 856
rect 125802 734 126278 856
rect 126446 734 126922 856
rect 127090 734 127566 856
rect 127734 734 128210 856
rect 128378 734 128854 856
rect 129022 734 129498 856
rect 129666 734 130142 856
rect 130310 734 130786 856
rect 130954 734 131430 856
rect 131598 734 131982 856
rect 132150 734 132626 856
rect 132794 734 133270 856
rect 133438 734 133914 856
rect 134082 734 134558 856
rect 134726 734 135202 856
rect 135370 734 135846 856
rect 136014 734 136490 856
rect 136658 734 137134 856
rect 137302 734 137778 856
rect 137946 734 138422 856
rect 138590 734 139066 856
rect 139234 734 139710 856
rect 139878 734 140262 856
rect 140430 734 140906 856
rect 141074 734 141550 856
rect 141718 734 142194 856
rect 142362 734 142838 856
rect 143006 734 143482 856
rect 143650 734 144126 856
rect 144294 734 144770 856
rect 144938 734 145414 856
rect 145582 734 146058 856
rect 146226 734 146702 856
rect 146870 734 147346 856
rect 147514 734 147990 856
rect 148158 734 148542 856
rect 148710 734 149186 856
rect 149354 734 149830 856
rect 149998 734 150474 856
rect 150642 734 151118 856
rect 151286 734 151762 856
rect 151930 734 152406 856
rect 152574 734 153050 856
rect 153218 734 153694 856
rect 153862 734 154338 856
rect 154506 734 154982 856
rect 155150 734 155626 856
rect 155794 734 156270 856
rect 156438 734 156822 856
rect 156990 734 157466 856
rect 157634 734 158110 856
rect 158278 734 158754 856
rect 158922 734 159398 856
rect 159566 734 160042 856
rect 160210 734 160686 856
rect 160854 734 161330 856
rect 161498 734 161974 856
rect 162142 734 162618 856
rect 162786 734 163262 856
rect 163430 734 163906 856
rect 164074 734 164458 856
rect 164626 734 165102 856
rect 165270 734 165746 856
rect 165914 734 166390 856
rect 166558 734 167034 856
rect 167202 734 167678 856
rect 167846 734 168322 856
rect 168490 734 168966 856
rect 169134 734 169610 856
rect 169778 734 170254 856
rect 170422 734 170898 856
rect 171066 734 171542 856
rect 171710 734 172186 856
rect 172354 734 172738 856
rect 172906 734 173382 856
rect 173550 734 174026 856
rect 174194 734 174670 856
rect 174838 734 175314 856
rect 175482 734 175958 856
rect 176126 734 176602 856
rect 176770 734 177246 856
rect 177414 734 177890 856
rect 178058 734 178534 856
rect 178702 734 179178 856
rect 179346 734 179822 856
rect 179990 734 180466 856
rect 180634 734 181018 856
rect 181186 734 181662 856
rect 181830 734 182306 856
rect 182474 734 182950 856
rect 183118 734 183594 856
rect 183762 734 184238 856
rect 184406 734 184882 856
rect 185050 734 185526 856
rect 185694 734 186170 856
rect 186338 734 186814 856
rect 186982 734 187458 856
rect 187626 734 188102 856
rect 188270 734 188746 856
rect 188914 734 189298 856
rect 189466 734 189942 856
rect 190110 734 190586 856
rect 190754 734 191230 856
rect 191398 734 191874 856
rect 192042 734 192518 856
rect 192686 734 193162 856
rect 193330 734 193806 856
rect 193974 734 194450 856
rect 194618 734 195094 856
rect 195262 734 195738 856
rect 195906 734 196382 856
rect 196550 734 197026 856
rect 197194 734 197578 856
rect 197746 734 198222 856
rect 198390 734 198866 856
rect 199034 734 199510 856
rect 199678 734 200154 856
rect 200322 734 200798 856
rect 200966 734 201442 856
rect 201610 734 202086 856
rect 202254 734 202730 856
rect 202898 734 203374 856
rect 203542 734 204018 856
rect 204186 734 204662 856
rect 204830 734 205306 856
rect 205474 734 205858 856
rect 206026 734 206502 856
rect 206670 734 207146 856
rect 207314 734 207790 856
rect 207958 734 208434 856
rect 208602 734 209078 856
rect 209246 734 209722 856
rect 209890 734 210366 856
rect 210534 734 211010 856
rect 211178 734 211654 856
rect 211822 734 212298 856
rect 212466 734 212942 856
rect 213110 734 213586 856
rect 213754 734 214138 856
rect 214306 734 214782 856
rect 214950 734 215426 856
rect 215594 734 216070 856
rect 216238 734 216714 856
rect 216882 734 217358 856
rect 217526 734 218002 856
rect 218170 734 218646 856
rect 218814 734 219290 856
rect 219458 734 219934 856
rect 220102 734 220578 856
rect 220746 734 221222 856
rect 221390 734 221866 856
rect 222034 734 222418 856
rect 222586 734 223062 856
rect 223230 734 223706 856
rect 223874 734 224350 856
rect 224518 734 224994 856
rect 225162 734 225638 856
rect 225806 734 226282 856
rect 226450 734 226926 856
rect 227094 734 227570 856
rect 227738 734 228214 856
rect 228382 734 228858 856
rect 229026 734 229502 856
rect 229670 734 230146 856
rect 230314 734 230698 856
rect 230866 734 231342 856
rect 231510 734 231986 856
rect 232154 734 232630 856
rect 232798 734 233274 856
rect 233442 734 233918 856
rect 234086 734 234562 856
rect 234730 734 235206 856
rect 235374 734 235850 856
rect 236018 734 236494 856
rect 236662 734 237138 856
rect 237306 734 237782 856
rect 237950 734 238334 856
rect 238502 734 238978 856
rect 239146 734 239622 856
rect 239790 734 240266 856
rect 240434 734 240910 856
rect 241078 734 241554 856
rect 241722 734 242198 856
rect 242366 734 242842 856
rect 243010 734 243486 856
rect 243654 734 244130 856
rect 244298 734 244774 856
rect 244942 734 245418 856
rect 245586 734 246062 856
rect 246230 734 246614 856
rect 246782 734 247258 856
rect 247426 734 247902 856
rect 248070 734 248546 856
rect 248714 734 249190 856
rect 249358 734 249834 856
rect 250002 734 250478 856
rect 250646 734 251122 856
rect 251290 734 251766 856
rect 251934 734 252410 856
rect 252578 734 253054 856
rect 253222 734 253698 856
rect 253866 734 254342 856
rect 254510 734 254894 856
rect 255062 734 255538 856
rect 255706 734 256182 856
rect 256350 734 256826 856
rect 256994 734 257470 856
rect 257638 734 258114 856
rect 258282 734 258758 856
rect 258926 734 259402 856
rect 259570 734 260046 856
rect 260214 734 260690 856
rect 260858 734 261334 856
rect 261502 734 261978 856
rect 262146 734 262622 856
rect 262790 734 263174 856
rect 263342 734 263818 856
rect 263986 734 264462 856
rect 264630 734 265106 856
rect 265274 734 265750 856
rect 265918 734 266394 856
rect 266562 734 267038 856
rect 267206 734 267682 856
rect 267850 734 268326 856
rect 268494 734 268970 856
rect 269138 734 269614 856
rect 269782 734 270258 856
rect 270426 734 270902 856
rect 271070 734 271454 856
rect 271622 734 272098 856
rect 272266 734 272742 856
rect 272910 734 273386 856
rect 273554 734 274030 856
rect 274198 734 274674 856
rect 274842 734 275318 856
rect 275486 734 275962 856
rect 276130 734 276606 856
rect 276774 734 277250 856
rect 277418 734 277894 856
rect 278062 734 278538 856
rect 278706 734 279182 856
rect 279350 734 279734 856
rect 279902 734 280378 856
rect 280546 734 281022 856
rect 281190 734 281666 856
rect 281834 734 282310 856
rect 282478 734 282954 856
rect 283122 734 283598 856
rect 283766 734 284242 856
rect 284410 734 284886 856
rect 285054 734 285530 856
rect 285698 734 286174 856
rect 286342 734 286818 856
rect 286986 734 287462 856
rect 287630 734 288014 856
rect 288182 734 288658 856
rect 288826 734 289302 856
rect 289470 734 289946 856
rect 290114 734 290590 856
rect 290758 734 291234 856
rect 291402 734 291878 856
rect 292046 734 292522 856
rect 292690 734 293166 856
rect 293334 734 293810 856
rect 293978 734 294454 856
rect 294622 734 295098 856
rect 295266 734 295742 856
rect 295910 734 296294 856
rect 296462 734 296938 856
rect 297106 734 297582 856
rect 297750 734 298226 856
rect 298394 734 298870 856
rect 299038 734 299514 856
rect 299682 734 300158 856
rect 300326 734 300802 856
rect 300970 734 301446 856
rect 301614 734 302090 856
rect 302258 734 302734 856
rect 302902 734 303378 856
rect 303546 734 304022 856
rect 304190 734 304574 856
rect 304742 734 305218 856
rect 305386 734 305862 856
rect 306030 734 306506 856
rect 306674 734 307150 856
rect 307318 734 307794 856
rect 307962 734 308438 856
rect 308606 734 309082 856
rect 309250 734 309726 856
rect 309894 734 310370 856
rect 310538 734 311014 856
<< obsm3 >>
rect 289 2143 296368 311745
<< metal4 >>
rect 4208 2128 4528 311760
rect 19568 2128 19888 311760
rect 34928 2128 35248 311760
rect 50288 2128 50608 311760
rect 65648 2128 65968 311760
rect 81008 2128 81328 311760
rect 96368 2128 96688 311760
rect 111728 2128 112048 311760
rect 127088 2128 127408 311760
rect 142448 2128 142768 311760
rect 157808 2128 158128 311760
rect 173168 2128 173488 311760
rect 188528 2128 188848 311760
rect 203888 2128 204208 311760
rect 219248 2128 219568 311760
rect 234608 2128 234928 311760
rect 249968 2128 250288 311760
rect 265328 2128 265648 311760
rect 280688 2128 281008 311760
rect 296048 2128 296368 311760
<< obsm4 >>
rect 18827 26827 19488 269381
rect 19968 26827 34848 269381
rect 35328 26827 50208 269381
rect 50688 26827 65568 269381
rect 66048 26827 80928 269381
rect 81408 26827 96288 269381
rect 96768 26827 111648 269381
rect 112128 26827 127008 269381
rect 127488 26827 142368 269381
rect 142848 26827 157728 269381
rect 158208 26827 173088 269381
rect 173568 26827 188448 269381
rect 188928 26827 203808 269381
rect 204288 26827 219168 269381
rect 219648 26827 234528 269381
rect 235008 26827 249888 269381
rect 250368 26827 265248 269381
rect 265728 26827 277045 269381
<< labels >>
rlabel metal2 s 1306 313367 1362 314167 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 83370 313367 83426 314167 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 91558 313367 91614 314167 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 99838 313367 99894 314167 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 108026 313367 108082 314167 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 116214 313367 116270 314167 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 124402 313367 124458 314167 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 132682 313367 132738 314167 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 140870 313367 140926 314167 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 149058 313367 149114 314167 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 157338 313367 157394 314167 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 9494 313367 9550 314167 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 165526 313367 165582 314167 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 173714 313367 173770 314167 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 181902 313367 181958 314167 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 190182 313367 190238 314167 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 198370 313367 198426 314167 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 206558 313367 206614 314167 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 214746 313367 214802 314167 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 223026 313367 223082 314167 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 231214 313367 231270 314167 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 239402 313367 239458 314167 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 17682 313367 17738 314167 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 247590 313367 247646 314167 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 255870 313367 255926 314167 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 264058 313367 264114 314167 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 272246 313367 272302 314167 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 280434 313367 280490 314167 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 288714 313367 288770 314167 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 296902 313367 296958 314167 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 305090 313367 305146 314167 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 25870 313367 25926 314167 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 34150 313367 34206 314167 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 42338 313367 42394 314167 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 50526 313367 50582 314167 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 58714 313367 58770 314167 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 66994 313367 67050 314167 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 75182 313367 75238 314167 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3974 313367 4030 314167 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 86130 313367 86186 314167 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 94318 313367 94374 314167 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 102506 313367 102562 314167 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 110786 313367 110842 314167 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 118974 313367 119030 314167 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 127162 313367 127218 314167 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 135350 313367 135406 314167 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 143630 313367 143686 314167 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 151818 313367 151874 314167 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 160006 313367 160062 314167 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 12254 313367 12310 314167 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 168286 313367 168342 314167 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 176474 313367 176530 314167 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 184662 313367 184718 314167 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 192850 313367 192906 314167 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 201130 313367 201186 314167 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 209318 313367 209374 314167 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 217506 313367 217562 314167 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 225694 313367 225750 314167 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 233974 313367 234030 314167 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 242162 313367 242218 314167 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 20442 313367 20498 314167 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 250350 313367 250406 314167 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 258538 313367 258594 314167 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 266818 313367 266874 314167 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 275006 313367 275062 314167 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 283194 313367 283250 314167 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 291382 313367 291438 314167 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 299662 313367 299718 314167 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 307850 313367 307906 314167 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 28630 313367 28686 314167 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 36818 313367 36874 314167 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 45098 313367 45154 314167 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 53286 313367 53342 314167 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 61474 313367 61530 314167 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 69662 313367 69718 314167 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 77942 313367 77998 314167 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 6734 313367 6790 314167 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 88890 313367 88946 314167 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 97078 313367 97134 314167 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 105266 313367 105322 314167 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 113454 313367 113510 314167 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 121734 313367 121790 314167 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 129922 313367 129978 314167 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 138110 313367 138166 314167 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 146298 313367 146354 314167 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 154578 313367 154634 314167 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 162766 313367 162822 314167 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 14922 313367 14978 314167 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 170954 313367 171010 314167 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 179234 313367 179290 314167 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 187422 313367 187478 314167 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 195610 313367 195666 314167 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 203798 313367 203854 314167 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 212078 313367 212134 314167 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 220266 313367 220322 314167 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 228454 313367 228510 314167 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 236642 313367 236698 314167 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 244922 313367 244978 314167 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 23202 313367 23258 314167 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 253110 313367 253166 314167 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 261298 313367 261354 314167 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 269486 313367 269542 314167 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 277766 313367 277822 314167 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 285954 313367 286010 314167 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 294142 313367 294198 314167 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 302330 313367 302386 314167 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 310610 313367 310666 314167 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 31390 313367 31446 314167 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 39578 313367 39634 314167 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 47766 313367 47822 314167 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 56046 313367 56102 314167 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 64234 313367 64290 314167 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 72422 313367 72478 314167 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 80610 313367 80666 314167 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 67730 0 67786 800 6 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 258814 0 258870 800 6 la_data_in[100]
port 116 nsew signal input
rlabel metal2 s 260746 0 260802 800 6 la_data_in[101]
port 117 nsew signal input
rlabel metal2 s 262678 0 262734 800 6 la_data_in[102]
port 118 nsew signal input
rlabel metal2 s 264518 0 264574 800 6 la_data_in[103]
port 119 nsew signal input
rlabel metal2 s 266450 0 266506 800 6 la_data_in[104]
port 120 nsew signal input
rlabel metal2 s 268382 0 268438 800 6 la_data_in[105]
port 121 nsew signal input
rlabel metal2 s 270314 0 270370 800 6 la_data_in[106]
port 122 nsew signal input
rlabel metal2 s 272154 0 272210 800 6 la_data_in[107]
port 123 nsew signal input
rlabel metal2 s 274086 0 274142 800 6 la_data_in[108]
port 124 nsew signal input
rlabel metal2 s 276018 0 276074 800 6 la_data_in[109]
port 125 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_data_in[10]
port 126 nsew signal input
rlabel metal2 s 277950 0 278006 800 6 la_data_in[110]
port 127 nsew signal input
rlabel metal2 s 279790 0 279846 800 6 la_data_in[111]
port 128 nsew signal input
rlabel metal2 s 281722 0 281778 800 6 la_data_in[112]
port 129 nsew signal input
rlabel metal2 s 283654 0 283710 800 6 la_data_in[113]
port 130 nsew signal input
rlabel metal2 s 285586 0 285642 800 6 la_data_in[114]
port 131 nsew signal input
rlabel metal2 s 287518 0 287574 800 6 la_data_in[115]
port 132 nsew signal input
rlabel metal2 s 289358 0 289414 800 6 la_data_in[116]
port 133 nsew signal input
rlabel metal2 s 291290 0 291346 800 6 la_data_in[117]
port 134 nsew signal input
rlabel metal2 s 293222 0 293278 800 6 la_data_in[118]
port 135 nsew signal input
rlabel metal2 s 295154 0 295210 800 6 la_data_in[119]
port 136 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_data_in[11]
port 137 nsew signal input
rlabel metal2 s 296994 0 297050 800 6 la_data_in[120]
port 138 nsew signal input
rlabel metal2 s 298926 0 298982 800 6 la_data_in[121]
port 139 nsew signal input
rlabel metal2 s 300858 0 300914 800 6 la_data_in[122]
port 140 nsew signal input
rlabel metal2 s 302790 0 302846 800 6 la_data_in[123]
port 141 nsew signal input
rlabel metal2 s 304630 0 304686 800 6 la_data_in[124]
port 142 nsew signal input
rlabel metal2 s 306562 0 306618 800 6 la_data_in[125]
port 143 nsew signal input
rlabel metal2 s 308494 0 308550 800 6 la_data_in[126]
port 144 nsew signal input
rlabel metal2 s 310426 0 310482 800 6 la_data_in[127]
port 145 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_data_in[12]
port 146 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_data_in[13]
port 147 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 la_data_in[14]
port 148 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_data_in[15]
port 149 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_data_in[16]
port 150 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 la_data_in[17]
port 151 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 la_data_in[18]
port 152 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 la_data_in[19]
port 153 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_data_in[1]
port 154 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 la_data_in[20]
port 155 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 la_data_in[21]
port 156 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 la_data_in[22]
port 157 nsew signal input
rlabel metal2 s 111706 0 111762 800 6 la_data_in[23]
port 158 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_data_in[24]
port 159 nsew signal input
rlabel metal2 s 115478 0 115534 800 6 la_data_in[25]
port 160 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 la_data_in[26]
port 161 nsew signal input
rlabel metal2 s 119342 0 119398 800 6 la_data_in[27]
port 162 nsew signal input
rlabel metal2 s 121274 0 121330 800 6 la_data_in[28]
port 163 nsew signal input
rlabel metal2 s 123206 0 123262 800 6 la_data_in[29]
port 164 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 la_data_in[2]
port 165 nsew signal input
rlabel metal2 s 125046 0 125102 800 6 la_data_in[30]
port 166 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_data_in[31]
port 167 nsew signal input
rlabel metal2 s 128910 0 128966 800 6 la_data_in[32]
port 168 nsew signal input
rlabel metal2 s 130842 0 130898 800 6 la_data_in[33]
port 169 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 la_data_in[34]
port 170 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 la_data_in[35]
port 171 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 la_data_in[36]
port 172 nsew signal input
rlabel metal2 s 138478 0 138534 800 6 la_data_in[37]
port 173 nsew signal input
rlabel metal2 s 140318 0 140374 800 6 la_data_in[38]
port 174 nsew signal input
rlabel metal2 s 142250 0 142306 800 6 la_data_in[39]
port 175 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 la_data_in[3]
port 176 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 la_data_in[40]
port 177 nsew signal input
rlabel metal2 s 146114 0 146170 800 6 la_data_in[41]
port 178 nsew signal input
rlabel metal2 s 148046 0 148102 800 6 la_data_in[42]
port 179 nsew signal input
rlabel metal2 s 149886 0 149942 800 6 la_data_in[43]
port 180 nsew signal input
rlabel metal2 s 151818 0 151874 800 6 la_data_in[44]
port 181 nsew signal input
rlabel metal2 s 153750 0 153806 800 6 la_data_in[45]
port 182 nsew signal input
rlabel metal2 s 155682 0 155738 800 6 la_data_in[46]
port 183 nsew signal input
rlabel metal2 s 157522 0 157578 800 6 la_data_in[47]
port 184 nsew signal input
rlabel metal2 s 159454 0 159510 800 6 la_data_in[48]
port 185 nsew signal input
rlabel metal2 s 161386 0 161442 800 6 la_data_in[49]
port 186 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_data_in[4]
port 187 nsew signal input
rlabel metal2 s 163318 0 163374 800 6 la_data_in[50]
port 188 nsew signal input
rlabel metal2 s 165158 0 165214 800 6 la_data_in[51]
port 189 nsew signal input
rlabel metal2 s 167090 0 167146 800 6 la_data_in[52]
port 190 nsew signal input
rlabel metal2 s 169022 0 169078 800 6 la_data_in[53]
port 191 nsew signal input
rlabel metal2 s 170954 0 171010 800 6 la_data_in[54]
port 192 nsew signal input
rlabel metal2 s 172794 0 172850 800 6 la_data_in[55]
port 193 nsew signal input
rlabel metal2 s 174726 0 174782 800 6 la_data_in[56]
port 194 nsew signal input
rlabel metal2 s 176658 0 176714 800 6 la_data_in[57]
port 195 nsew signal input
rlabel metal2 s 178590 0 178646 800 6 la_data_in[58]
port 196 nsew signal input
rlabel metal2 s 180522 0 180578 800 6 la_data_in[59]
port 197 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 la_data_in[5]
port 198 nsew signal input
rlabel metal2 s 182362 0 182418 800 6 la_data_in[60]
port 199 nsew signal input
rlabel metal2 s 184294 0 184350 800 6 la_data_in[61]
port 200 nsew signal input
rlabel metal2 s 186226 0 186282 800 6 la_data_in[62]
port 201 nsew signal input
rlabel metal2 s 188158 0 188214 800 6 la_data_in[63]
port 202 nsew signal input
rlabel metal2 s 189998 0 190054 800 6 la_data_in[64]
port 203 nsew signal input
rlabel metal2 s 191930 0 191986 800 6 la_data_in[65]
port 204 nsew signal input
rlabel metal2 s 193862 0 193918 800 6 la_data_in[66]
port 205 nsew signal input
rlabel metal2 s 195794 0 195850 800 6 la_data_in[67]
port 206 nsew signal input
rlabel metal2 s 197634 0 197690 800 6 la_data_in[68]
port 207 nsew signal input
rlabel metal2 s 199566 0 199622 800 6 la_data_in[69]
port 208 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_data_in[6]
port 209 nsew signal input
rlabel metal2 s 201498 0 201554 800 6 la_data_in[70]
port 210 nsew signal input
rlabel metal2 s 203430 0 203486 800 6 la_data_in[71]
port 211 nsew signal input
rlabel metal2 s 205362 0 205418 800 6 la_data_in[72]
port 212 nsew signal input
rlabel metal2 s 207202 0 207258 800 6 la_data_in[73]
port 213 nsew signal input
rlabel metal2 s 209134 0 209190 800 6 la_data_in[74]
port 214 nsew signal input
rlabel metal2 s 211066 0 211122 800 6 la_data_in[75]
port 215 nsew signal input
rlabel metal2 s 212998 0 213054 800 6 la_data_in[76]
port 216 nsew signal input
rlabel metal2 s 214838 0 214894 800 6 la_data_in[77]
port 217 nsew signal input
rlabel metal2 s 216770 0 216826 800 6 la_data_in[78]
port 218 nsew signal input
rlabel metal2 s 218702 0 218758 800 6 la_data_in[79]
port 219 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_data_in[7]
port 220 nsew signal input
rlabel metal2 s 220634 0 220690 800 6 la_data_in[80]
port 221 nsew signal input
rlabel metal2 s 222474 0 222530 800 6 la_data_in[81]
port 222 nsew signal input
rlabel metal2 s 224406 0 224462 800 6 la_data_in[82]
port 223 nsew signal input
rlabel metal2 s 226338 0 226394 800 6 la_data_in[83]
port 224 nsew signal input
rlabel metal2 s 228270 0 228326 800 6 la_data_in[84]
port 225 nsew signal input
rlabel metal2 s 230202 0 230258 800 6 la_data_in[85]
port 226 nsew signal input
rlabel metal2 s 232042 0 232098 800 6 la_data_in[86]
port 227 nsew signal input
rlabel metal2 s 233974 0 234030 800 6 la_data_in[87]
port 228 nsew signal input
rlabel metal2 s 235906 0 235962 800 6 la_data_in[88]
port 229 nsew signal input
rlabel metal2 s 237838 0 237894 800 6 la_data_in[89]
port 230 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 la_data_in[8]
port 231 nsew signal input
rlabel metal2 s 239678 0 239734 800 6 la_data_in[90]
port 232 nsew signal input
rlabel metal2 s 241610 0 241666 800 6 la_data_in[91]
port 233 nsew signal input
rlabel metal2 s 243542 0 243598 800 6 la_data_in[92]
port 234 nsew signal input
rlabel metal2 s 245474 0 245530 800 6 la_data_in[93]
port 235 nsew signal input
rlabel metal2 s 247314 0 247370 800 6 la_data_in[94]
port 236 nsew signal input
rlabel metal2 s 249246 0 249302 800 6 la_data_in[95]
port 237 nsew signal input
rlabel metal2 s 251178 0 251234 800 6 la_data_in[96]
port 238 nsew signal input
rlabel metal2 s 253110 0 253166 800 6 la_data_in[97]
port 239 nsew signal input
rlabel metal2 s 254950 0 255006 800 6 la_data_in[98]
port 240 nsew signal input
rlabel metal2 s 256882 0 256938 800 6 la_data_in[99]
port 241 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_data_in[9]
port 242 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_data_out[0]
port 243 nsew signal output
rlabel metal2 s 259458 0 259514 800 6 la_data_out[100]
port 244 nsew signal output
rlabel metal2 s 261390 0 261446 800 6 la_data_out[101]
port 245 nsew signal output
rlabel metal2 s 263230 0 263286 800 6 la_data_out[102]
port 246 nsew signal output
rlabel metal2 s 265162 0 265218 800 6 la_data_out[103]
port 247 nsew signal output
rlabel metal2 s 267094 0 267150 800 6 la_data_out[104]
port 248 nsew signal output
rlabel metal2 s 269026 0 269082 800 6 la_data_out[105]
port 249 nsew signal output
rlabel metal2 s 270958 0 271014 800 6 la_data_out[106]
port 250 nsew signal output
rlabel metal2 s 272798 0 272854 800 6 la_data_out[107]
port 251 nsew signal output
rlabel metal2 s 274730 0 274786 800 6 la_data_out[108]
port 252 nsew signal output
rlabel metal2 s 276662 0 276718 800 6 la_data_out[109]
port 253 nsew signal output
rlabel metal2 s 87510 0 87566 800 6 la_data_out[10]
port 254 nsew signal output
rlabel metal2 s 278594 0 278650 800 6 la_data_out[110]
port 255 nsew signal output
rlabel metal2 s 280434 0 280490 800 6 la_data_out[111]
port 256 nsew signal output
rlabel metal2 s 282366 0 282422 800 6 la_data_out[112]
port 257 nsew signal output
rlabel metal2 s 284298 0 284354 800 6 la_data_out[113]
port 258 nsew signal output
rlabel metal2 s 286230 0 286286 800 6 la_data_out[114]
port 259 nsew signal output
rlabel metal2 s 288070 0 288126 800 6 la_data_out[115]
port 260 nsew signal output
rlabel metal2 s 290002 0 290058 800 6 la_data_out[116]
port 261 nsew signal output
rlabel metal2 s 291934 0 291990 800 6 la_data_out[117]
port 262 nsew signal output
rlabel metal2 s 293866 0 293922 800 6 la_data_out[118]
port 263 nsew signal output
rlabel metal2 s 295798 0 295854 800 6 la_data_out[119]
port 264 nsew signal output
rlabel metal2 s 89442 0 89498 800 6 la_data_out[11]
port 265 nsew signal output
rlabel metal2 s 297638 0 297694 800 6 la_data_out[120]
port 266 nsew signal output
rlabel metal2 s 299570 0 299626 800 6 la_data_out[121]
port 267 nsew signal output
rlabel metal2 s 301502 0 301558 800 6 la_data_out[122]
port 268 nsew signal output
rlabel metal2 s 303434 0 303490 800 6 la_data_out[123]
port 269 nsew signal output
rlabel metal2 s 305274 0 305330 800 6 la_data_out[124]
port 270 nsew signal output
rlabel metal2 s 307206 0 307262 800 6 la_data_out[125]
port 271 nsew signal output
rlabel metal2 s 309138 0 309194 800 6 la_data_out[126]
port 272 nsew signal output
rlabel metal2 s 311070 0 311126 800 6 la_data_out[127]
port 273 nsew signal output
rlabel metal2 s 91282 0 91338 800 6 la_data_out[12]
port 274 nsew signal output
rlabel metal2 s 93214 0 93270 800 6 la_data_out[13]
port 275 nsew signal output
rlabel metal2 s 95146 0 95202 800 6 la_data_out[14]
port 276 nsew signal output
rlabel metal2 s 97078 0 97134 800 6 la_data_out[15]
port 277 nsew signal output
rlabel metal2 s 98918 0 98974 800 6 la_data_out[16]
port 278 nsew signal output
rlabel metal2 s 100850 0 100906 800 6 la_data_out[17]
port 279 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 la_data_out[18]
port 280 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 la_data_out[19]
port 281 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 la_data_out[1]
port 282 nsew signal output
rlabel metal2 s 106646 0 106702 800 6 la_data_out[20]
port 283 nsew signal output
rlabel metal2 s 108486 0 108542 800 6 la_data_out[21]
port 284 nsew signal output
rlabel metal2 s 110418 0 110474 800 6 la_data_out[22]
port 285 nsew signal output
rlabel metal2 s 112350 0 112406 800 6 la_data_out[23]
port 286 nsew signal output
rlabel metal2 s 114282 0 114338 800 6 la_data_out[24]
port 287 nsew signal output
rlabel metal2 s 116122 0 116178 800 6 la_data_out[25]
port 288 nsew signal output
rlabel metal2 s 118054 0 118110 800 6 la_data_out[26]
port 289 nsew signal output
rlabel metal2 s 119986 0 120042 800 6 la_data_out[27]
port 290 nsew signal output
rlabel metal2 s 121918 0 121974 800 6 la_data_out[28]
port 291 nsew signal output
rlabel metal2 s 123758 0 123814 800 6 la_data_out[29]
port 292 nsew signal output
rlabel metal2 s 72238 0 72294 800 6 la_data_out[2]
port 293 nsew signal output
rlabel metal2 s 125690 0 125746 800 6 la_data_out[30]
port 294 nsew signal output
rlabel metal2 s 127622 0 127678 800 6 la_data_out[31]
port 295 nsew signal output
rlabel metal2 s 129554 0 129610 800 6 la_data_out[32]
port 296 nsew signal output
rlabel metal2 s 131486 0 131542 800 6 la_data_out[33]
port 297 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 la_data_out[34]
port 298 nsew signal output
rlabel metal2 s 135258 0 135314 800 6 la_data_out[35]
port 299 nsew signal output
rlabel metal2 s 137190 0 137246 800 6 la_data_out[36]
port 300 nsew signal output
rlabel metal2 s 139122 0 139178 800 6 la_data_out[37]
port 301 nsew signal output
rlabel metal2 s 140962 0 141018 800 6 la_data_out[38]
port 302 nsew signal output
rlabel metal2 s 142894 0 142950 800 6 la_data_out[39]
port 303 nsew signal output
rlabel metal2 s 74170 0 74226 800 6 la_data_out[3]
port 304 nsew signal output
rlabel metal2 s 144826 0 144882 800 6 la_data_out[40]
port 305 nsew signal output
rlabel metal2 s 146758 0 146814 800 6 la_data_out[41]
port 306 nsew signal output
rlabel metal2 s 148598 0 148654 800 6 la_data_out[42]
port 307 nsew signal output
rlabel metal2 s 150530 0 150586 800 6 la_data_out[43]
port 308 nsew signal output
rlabel metal2 s 152462 0 152518 800 6 la_data_out[44]
port 309 nsew signal output
rlabel metal2 s 154394 0 154450 800 6 la_data_out[45]
port 310 nsew signal output
rlabel metal2 s 156326 0 156382 800 6 la_data_out[46]
port 311 nsew signal output
rlabel metal2 s 158166 0 158222 800 6 la_data_out[47]
port 312 nsew signal output
rlabel metal2 s 160098 0 160154 800 6 la_data_out[48]
port 313 nsew signal output
rlabel metal2 s 162030 0 162086 800 6 la_data_out[49]
port 314 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 la_data_out[4]
port 315 nsew signal output
rlabel metal2 s 163962 0 164018 800 6 la_data_out[50]
port 316 nsew signal output
rlabel metal2 s 165802 0 165858 800 6 la_data_out[51]
port 317 nsew signal output
rlabel metal2 s 167734 0 167790 800 6 la_data_out[52]
port 318 nsew signal output
rlabel metal2 s 169666 0 169722 800 6 la_data_out[53]
port 319 nsew signal output
rlabel metal2 s 171598 0 171654 800 6 la_data_out[54]
port 320 nsew signal output
rlabel metal2 s 173438 0 173494 800 6 la_data_out[55]
port 321 nsew signal output
rlabel metal2 s 175370 0 175426 800 6 la_data_out[56]
port 322 nsew signal output
rlabel metal2 s 177302 0 177358 800 6 la_data_out[57]
port 323 nsew signal output
rlabel metal2 s 179234 0 179290 800 6 la_data_out[58]
port 324 nsew signal output
rlabel metal2 s 181074 0 181130 800 6 la_data_out[59]
port 325 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 la_data_out[5]
port 326 nsew signal output
rlabel metal2 s 183006 0 183062 800 6 la_data_out[60]
port 327 nsew signal output
rlabel metal2 s 184938 0 184994 800 6 la_data_out[61]
port 328 nsew signal output
rlabel metal2 s 186870 0 186926 800 6 la_data_out[62]
port 329 nsew signal output
rlabel metal2 s 188802 0 188858 800 6 la_data_out[63]
port 330 nsew signal output
rlabel metal2 s 190642 0 190698 800 6 la_data_out[64]
port 331 nsew signal output
rlabel metal2 s 192574 0 192630 800 6 la_data_out[65]
port 332 nsew signal output
rlabel metal2 s 194506 0 194562 800 6 la_data_out[66]
port 333 nsew signal output
rlabel metal2 s 196438 0 196494 800 6 la_data_out[67]
port 334 nsew signal output
rlabel metal2 s 198278 0 198334 800 6 la_data_out[68]
port 335 nsew signal output
rlabel metal2 s 200210 0 200266 800 6 la_data_out[69]
port 336 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 la_data_out[6]
port 337 nsew signal output
rlabel metal2 s 202142 0 202198 800 6 la_data_out[70]
port 338 nsew signal output
rlabel metal2 s 204074 0 204130 800 6 la_data_out[71]
port 339 nsew signal output
rlabel metal2 s 205914 0 205970 800 6 la_data_out[72]
port 340 nsew signal output
rlabel metal2 s 207846 0 207902 800 6 la_data_out[73]
port 341 nsew signal output
rlabel metal2 s 209778 0 209834 800 6 la_data_out[74]
port 342 nsew signal output
rlabel metal2 s 211710 0 211766 800 6 la_data_out[75]
port 343 nsew signal output
rlabel metal2 s 213642 0 213698 800 6 la_data_out[76]
port 344 nsew signal output
rlabel metal2 s 215482 0 215538 800 6 la_data_out[77]
port 345 nsew signal output
rlabel metal2 s 217414 0 217470 800 6 la_data_out[78]
port 346 nsew signal output
rlabel metal2 s 219346 0 219402 800 6 la_data_out[79]
port 347 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 la_data_out[7]
port 348 nsew signal output
rlabel metal2 s 221278 0 221334 800 6 la_data_out[80]
port 349 nsew signal output
rlabel metal2 s 223118 0 223174 800 6 la_data_out[81]
port 350 nsew signal output
rlabel metal2 s 225050 0 225106 800 6 la_data_out[82]
port 351 nsew signal output
rlabel metal2 s 226982 0 227038 800 6 la_data_out[83]
port 352 nsew signal output
rlabel metal2 s 228914 0 228970 800 6 la_data_out[84]
port 353 nsew signal output
rlabel metal2 s 230754 0 230810 800 6 la_data_out[85]
port 354 nsew signal output
rlabel metal2 s 232686 0 232742 800 6 la_data_out[86]
port 355 nsew signal output
rlabel metal2 s 234618 0 234674 800 6 la_data_out[87]
port 356 nsew signal output
rlabel metal2 s 236550 0 236606 800 6 la_data_out[88]
port 357 nsew signal output
rlabel metal2 s 238390 0 238446 800 6 la_data_out[89]
port 358 nsew signal output
rlabel metal2 s 83646 0 83702 800 6 la_data_out[8]
port 359 nsew signal output
rlabel metal2 s 240322 0 240378 800 6 la_data_out[90]
port 360 nsew signal output
rlabel metal2 s 242254 0 242310 800 6 la_data_out[91]
port 361 nsew signal output
rlabel metal2 s 244186 0 244242 800 6 la_data_out[92]
port 362 nsew signal output
rlabel metal2 s 246118 0 246174 800 6 la_data_out[93]
port 363 nsew signal output
rlabel metal2 s 247958 0 248014 800 6 la_data_out[94]
port 364 nsew signal output
rlabel metal2 s 249890 0 249946 800 6 la_data_out[95]
port 365 nsew signal output
rlabel metal2 s 251822 0 251878 800 6 la_data_out[96]
port 366 nsew signal output
rlabel metal2 s 253754 0 253810 800 6 la_data_out[97]
port 367 nsew signal output
rlabel metal2 s 255594 0 255650 800 6 la_data_out[98]
port 368 nsew signal output
rlabel metal2 s 257526 0 257582 800 6 la_data_out[99]
port 369 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 la_data_out[9]
port 370 nsew signal output
rlabel metal2 s 69018 0 69074 800 6 la_oen[0]
port 371 nsew signal input
rlabel metal2 s 260102 0 260158 800 6 la_oen[100]
port 372 nsew signal input
rlabel metal2 s 262034 0 262090 800 6 la_oen[101]
port 373 nsew signal input
rlabel metal2 s 263874 0 263930 800 6 la_oen[102]
port 374 nsew signal input
rlabel metal2 s 265806 0 265862 800 6 la_oen[103]
port 375 nsew signal input
rlabel metal2 s 267738 0 267794 800 6 la_oen[104]
port 376 nsew signal input
rlabel metal2 s 269670 0 269726 800 6 la_oen[105]
port 377 nsew signal input
rlabel metal2 s 271510 0 271566 800 6 la_oen[106]
port 378 nsew signal input
rlabel metal2 s 273442 0 273498 800 6 la_oen[107]
port 379 nsew signal input
rlabel metal2 s 275374 0 275430 800 6 la_oen[108]
port 380 nsew signal input
rlabel metal2 s 277306 0 277362 800 6 la_oen[109]
port 381 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 la_oen[10]
port 382 nsew signal input
rlabel metal2 s 279238 0 279294 800 6 la_oen[110]
port 383 nsew signal input
rlabel metal2 s 281078 0 281134 800 6 la_oen[111]
port 384 nsew signal input
rlabel metal2 s 283010 0 283066 800 6 la_oen[112]
port 385 nsew signal input
rlabel metal2 s 284942 0 284998 800 6 la_oen[113]
port 386 nsew signal input
rlabel metal2 s 286874 0 286930 800 6 la_oen[114]
port 387 nsew signal input
rlabel metal2 s 288714 0 288770 800 6 la_oen[115]
port 388 nsew signal input
rlabel metal2 s 290646 0 290702 800 6 la_oen[116]
port 389 nsew signal input
rlabel metal2 s 292578 0 292634 800 6 la_oen[117]
port 390 nsew signal input
rlabel metal2 s 294510 0 294566 800 6 la_oen[118]
port 391 nsew signal input
rlabel metal2 s 296350 0 296406 800 6 la_oen[119]
port 392 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_oen[11]
port 393 nsew signal input
rlabel metal2 s 298282 0 298338 800 6 la_oen[120]
port 394 nsew signal input
rlabel metal2 s 300214 0 300270 800 6 la_oen[121]
port 395 nsew signal input
rlabel metal2 s 302146 0 302202 800 6 la_oen[122]
port 396 nsew signal input
rlabel metal2 s 304078 0 304134 800 6 la_oen[123]
port 397 nsew signal input
rlabel metal2 s 305918 0 305974 800 6 la_oen[124]
port 398 nsew signal input
rlabel metal2 s 307850 0 307906 800 6 la_oen[125]
port 399 nsew signal input
rlabel metal2 s 309782 0 309838 800 6 la_oen[126]
port 400 nsew signal input
rlabel metal2 s 311714 0 311770 800 6 la_oen[127]
port 401 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_oen[12]
port 402 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_oen[13]
port 403 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_oen[14]
port 404 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 la_oen[15]
port 405 nsew signal input
rlabel metal2 s 99562 0 99618 800 6 la_oen[16]
port 406 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 la_oen[17]
port 407 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 la_oen[18]
port 408 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 la_oen[19]
port 409 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_oen[1]
port 410 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 la_oen[20]
port 411 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_oen[21]
port 412 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 la_oen[22]
port 413 nsew signal input
rlabel metal2 s 112994 0 113050 800 6 la_oen[23]
port 414 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 la_oen[24]
port 415 nsew signal input
rlabel metal2 s 116766 0 116822 800 6 la_oen[25]
port 416 nsew signal input
rlabel metal2 s 118698 0 118754 800 6 la_oen[26]
port 417 nsew signal input
rlabel metal2 s 120630 0 120686 800 6 la_oen[27]
port 418 nsew signal input
rlabel metal2 s 122562 0 122618 800 6 la_oen[28]
port 419 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 la_oen[29]
port 420 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 la_oen[2]
port 421 nsew signal input
rlabel metal2 s 126334 0 126390 800 6 la_oen[30]
port 422 nsew signal input
rlabel metal2 s 128266 0 128322 800 6 la_oen[31]
port 423 nsew signal input
rlabel metal2 s 130198 0 130254 800 6 la_oen[32]
port 424 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 la_oen[33]
port 425 nsew signal input
rlabel metal2 s 133970 0 134026 800 6 la_oen[34]
port 426 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 la_oen[35]
port 427 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 la_oen[36]
port 428 nsew signal input
rlabel metal2 s 139766 0 139822 800 6 la_oen[37]
port 429 nsew signal input
rlabel metal2 s 141606 0 141662 800 6 la_oen[38]
port 430 nsew signal input
rlabel metal2 s 143538 0 143594 800 6 la_oen[39]
port 431 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 la_oen[3]
port 432 nsew signal input
rlabel metal2 s 145470 0 145526 800 6 la_oen[40]
port 433 nsew signal input
rlabel metal2 s 147402 0 147458 800 6 la_oen[41]
port 434 nsew signal input
rlabel metal2 s 149242 0 149298 800 6 la_oen[42]
port 435 nsew signal input
rlabel metal2 s 151174 0 151230 800 6 la_oen[43]
port 436 nsew signal input
rlabel metal2 s 153106 0 153162 800 6 la_oen[44]
port 437 nsew signal input
rlabel metal2 s 155038 0 155094 800 6 la_oen[45]
port 438 nsew signal input
rlabel metal2 s 156878 0 156934 800 6 la_oen[46]
port 439 nsew signal input
rlabel metal2 s 158810 0 158866 800 6 la_oen[47]
port 440 nsew signal input
rlabel metal2 s 160742 0 160798 800 6 la_oen[48]
port 441 nsew signal input
rlabel metal2 s 162674 0 162730 800 6 la_oen[49]
port 442 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 la_oen[4]
port 443 nsew signal input
rlabel metal2 s 164514 0 164570 800 6 la_oen[50]
port 444 nsew signal input
rlabel metal2 s 166446 0 166502 800 6 la_oen[51]
port 445 nsew signal input
rlabel metal2 s 168378 0 168434 800 6 la_oen[52]
port 446 nsew signal input
rlabel metal2 s 170310 0 170366 800 6 la_oen[53]
port 447 nsew signal input
rlabel metal2 s 172242 0 172298 800 6 la_oen[54]
port 448 nsew signal input
rlabel metal2 s 174082 0 174138 800 6 la_oen[55]
port 449 nsew signal input
rlabel metal2 s 176014 0 176070 800 6 la_oen[56]
port 450 nsew signal input
rlabel metal2 s 177946 0 178002 800 6 la_oen[57]
port 451 nsew signal input
rlabel metal2 s 179878 0 179934 800 6 la_oen[58]
port 452 nsew signal input
rlabel metal2 s 181718 0 181774 800 6 la_oen[59]
port 453 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 la_oen[5]
port 454 nsew signal input
rlabel metal2 s 183650 0 183706 800 6 la_oen[60]
port 455 nsew signal input
rlabel metal2 s 185582 0 185638 800 6 la_oen[61]
port 456 nsew signal input
rlabel metal2 s 187514 0 187570 800 6 la_oen[62]
port 457 nsew signal input
rlabel metal2 s 189354 0 189410 800 6 la_oen[63]
port 458 nsew signal input
rlabel metal2 s 191286 0 191342 800 6 la_oen[64]
port 459 nsew signal input
rlabel metal2 s 193218 0 193274 800 6 la_oen[65]
port 460 nsew signal input
rlabel metal2 s 195150 0 195206 800 6 la_oen[66]
port 461 nsew signal input
rlabel metal2 s 197082 0 197138 800 6 la_oen[67]
port 462 nsew signal input
rlabel metal2 s 198922 0 198978 800 6 la_oen[68]
port 463 nsew signal input
rlabel metal2 s 200854 0 200910 800 6 la_oen[69]
port 464 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_oen[6]
port 465 nsew signal input
rlabel metal2 s 202786 0 202842 800 6 la_oen[70]
port 466 nsew signal input
rlabel metal2 s 204718 0 204774 800 6 la_oen[71]
port 467 nsew signal input
rlabel metal2 s 206558 0 206614 800 6 la_oen[72]
port 468 nsew signal input
rlabel metal2 s 208490 0 208546 800 6 la_oen[73]
port 469 nsew signal input
rlabel metal2 s 210422 0 210478 800 6 la_oen[74]
port 470 nsew signal input
rlabel metal2 s 212354 0 212410 800 6 la_oen[75]
port 471 nsew signal input
rlabel metal2 s 214194 0 214250 800 6 la_oen[76]
port 472 nsew signal input
rlabel metal2 s 216126 0 216182 800 6 la_oen[77]
port 473 nsew signal input
rlabel metal2 s 218058 0 218114 800 6 la_oen[78]
port 474 nsew signal input
rlabel metal2 s 219990 0 220046 800 6 la_oen[79]
port 475 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_oen[7]
port 476 nsew signal input
rlabel metal2 s 221922 0 221978 800 6 la_oen[80]
port 477 nsew signal input
rlabel metal2 s 223762 0 223818 800 6 la_oen[81]
port 478 nsew signal input
rlabel metal2 s 225694 0 225750 800 6 la_oen[82]
port 479 nsew signal input
rlabel metal2 s 227626 0 227682 800 6 la_oen[83]
port 480 nsew signal input
rlabel metal2 s 229558 0 229614 800 6 la_oen[84]
port 481 nsew signal input
rlabel metal2 s 231398 0 231454 800 6 la_oen[85]
port 482 nsew signal input
rlabel metal2 s 233330 0 233386 800 6 la_oen[86]
port 483 nsew signal input
rlabel metal2 s 235262 0 235318 800 6 la_oen[87]
port 484 nsew signal input
rlabel metal2 s 237194 0 237250 800 6 la_oen[88]
port 485 nsew signal input
rlabel metal2 s 239034 0 239090 800 6 la_oen[89]
port 486 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_oen[8]
port 487 nsew signal input
rlabel metal2 s 240966 0 241022 800 6 la_oen[90]
port 488 nsew signal input
rlabel metal2 s 242898 0 242954 800 6 la_oen[91]
port 489 nsew signal input
rlabel metal2 s 244830 0 244886 800 6 la_oen[92]
port 490 nsew signal input
rlabel metal2 s 246670 0 246726 800 6 la_oen[93]
port 491 nsew signal input
rlabel metal2 s 248602 0 248658 800 6 la_oen[94]
port 492 nsew signal input
rlabel metal2 s 250534 0 250590 800 6 la_oen[95]
port 493 nsew signal input
rlabel metal2 s 252466 0 252522 800 6 la_oen[96]
port 494 nsew signal input
rlabel metal2 s 254398 0 254454 800 6 la_oen[97]
port 495 nsew signal input
rlabel metal2 s 256238 0 256294 800 6 la_oen[98]
port 496 nsew signal input
rlabel metal2 s 258170 0 258226 800 6 la_oen[99]
port 497 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_oen[9]
port 498 nsew signal input
rlabel metal4 s 4208 2128 4528 311760 6 vccd1
port 499 nsew power input
rlabel metal4 s 34928 2128 35248 311760 6 vccd1
port 499 nsew power input
rlabel metal4 s 65648 2128 65968 311760 6 vccd1
port 499 nsew power input
rlabel metal4 s 96368 2128 96688 311760 6 vccd1
port 499 nsew power input
rlabel metal4 s 127088 2128 127408 311760 6 vccd1
port 499 nsew power input
rlabel metal4 s 157808 2128 158128 311760 6 vccd1
port 499 nsew power input
rlabel metal4 s 188528 2128 188848 311760 6 vccd1
port 499 nsew power input
rlabel metal4 s 219248 2128 219568 311760 6 vccd1
port 499 nsew power input
rlabel metal4 s 249968 2128 250288 311760 6 vccd1
port 499 nsew power input
rlabel metal4 s 280688 2128 281008 311760 6 vccd1
port 499 nsew power input
rlabel metal4 s 19568 2128 19888 311760 6 vssd1
port 500 nsew ground input
rlabel metal4 s 50288 2128 50608 311760 6 vssd1
port 500 nsew ground input
rlabel metal4 s 81008 2128 81328 311760 6 vssd1
port 500 nsew ground input
rlabel metal4 s 111728 2128 112048 311760 6 vssd1
port 500 nsew ground input
rlabel metal4 s 142448 2128 142768 311760 6 vssd1
port 500 nsew ground input
rlabel metal4 s 173168 2128 173488 311760 6 vssd1
port 500 nsew ground input
rlabel metal4 s 203888 2128 204208 311760 6 vssd1
port 500 nsew ground input
rlabel metal4 s 234608 2128 234928 311760 6 vssd1
port 500 nsew ground input
rlabel metal4 s 265328 2128 265648 311760 6 vssd1
port 500 nsew ground input
rlabel metal4 s 296048 2128 296368 311760 6 vssd1
port 500 nsew ground input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 501 nsew signal input
rlabel metal2 s 846 0 902 800 6 wb_rst_i
port 502 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_ack_o
port 503 nsew signal output
rlabel metal2 s 4066 0 4122 800 6 wbs_adr_i[0]
port 504 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 wbs_adr_i[10]
port 505 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 wbs_adr_i[11]
port 506 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 wbs_adr_i[12]
port 507 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 wbs_adr_i[13]
port 508 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wbs_adr_i[14]
port 509 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 wbs_adr_i[15]
port 510 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wbs_adr_i[16]
port 511 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 wbs_adr_i[17]
port 512 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 wbs_adr_i[18]
port 513 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 wbs_adr_i[19]
port 514 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_adr_i[1]
port 515 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 wbs_adr_i[20]
port 516 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 wbs_adr_i[21]
port 517 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 wbs_adr_i[22]
port 518 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 wbs_adr_i[23]
port 519 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 wbs_adr_i[24]
port 520 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 wbs_adr_i[25]
port 521 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 wbs_adr_i[26]
port 522 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 wbs_adr_i[27]
port 523 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 wbs_adr_i[28]
port 524 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 wbs_adr_i[29]
port 525 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_adr_i[2]
port 526 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 wbs_adr_i[30]
port 527 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 wbs_adr_i[31]
port 528 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wbs_adr_i[3]
port 529 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_adr_i[4]
port 530 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 wbs_adr_i[5]
port 531 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_adr_i[6]
port 532 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_adr_i[7]
port 533 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wbs_adr_i[8]
port 534 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 wbs_adr_i[9]
port 535 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_cyc_i
port 536 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_i[0]
port 537 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_dat_i[10]
port 538 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 wbs_dat_i[11]
port 539 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_i[12]
port 540 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_i[13]
port 541 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 wbs_dat_i[14]
port 542 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_dat_i[15]
port 543 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_dat_i[16]
port 544 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 wbs_dat_i[17]
port 545 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 wbs_dat_i[18]
port 546 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 wbs_dat_i[19]
port 547 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 wbs_dat_i[1]
port 548 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 wbs_dat_i[20]
port 549 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 wbs_dat_i[21]
port 550 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 wbs_dat_i[22]
port 551 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 wbs_dat_i[23]
port 552 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 wbs_dat_i[24]
port 553 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 wbs_dat_i[25]
port 554 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 wbs_dat_i[26]
port 555 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 wbs_dat_i[27]
port 556 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 wbs_dat_i[28]
port 557 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 wbs_dat_i[29]
port 558 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_i[2]
port 559 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 wbs_dat_i[30]
port 560 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 wbs_dat_i[31]
port 561 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_i[3]
port 562 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_dat_i[4]
port 563 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_dat_i[5]
port 564 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_i[6]
port 565 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_i[7]
port 566 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_i[8]
port 567 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_dat_i[9]
port 568 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_o[0]
port 569 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_o[10]
port 570 nsew signal output
rlabel metal2 s 28906 0 28962 800 6 wbs_dat_o[11]
port 571 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 wbs_dat_o[12]
port 572 nsew signal output
rlabel metal2 s 32770 0 32826 800 6 wbs_dat_o[13]
port 573 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 wbs_dat_o[14]
port 574 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 wbs_dat_o[15]
port 575 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 wbs_dat_o[16]
port 576 nsew signal output
rlabel metal2 s 40406 0 40462 800 6 wbs_dat_o[17]
port 577 nsew signal output
rlabel metal2 s 42246 0 42302 800 6 wbs_dat_o[18]
port 578 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 wbs_dat_o[19]
port 579 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_o[1]
port 580 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 wbs_dat_o[20]
port 581 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 wbs_dat_o[21]
port 582 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 wbs_dat_o[22]
port 583 nsew signal output
rlabel metal2 s 51814 0 51870 800 6 wbs_dat_o[23]
port 584 nsew signal output
rlabel metal2 s 53746 0 53802 800 6 wbs_dat_o[24]
port 585 nsew signal output
rlabel metal2 s 55678 0 55734 800 6 wbs_dat_o[25]
port 586 nsew signal output
rlabel metal2 s 57610 0 57666 800 6 wbs_dat_o[26]
port 587 nsew signal output
rlabel metal2 s 59450 0 59506 800 6 wbs_dat_o[27]
port 588 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 wbs_dat_o[28]
port 589 nsew signal output
rlabel metal2 s 63314 0 63370 800 6 wbs_dat_o[29]
port 590 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_o[2]
port 591 nsew signal output
rlabel metal2 s 65246 0 65302 800 6 wbs_dat_o[30]
port 592 nsew signal output
rlabel metal2 s 67086 0 67142 800 6 wbs_dat_o[31]
port 593 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_o[3]
port 594 nsew signal output
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_o[4]
port 595 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_o[5]
port 596 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_o[6]
port 597 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 wbs_dat_o[7]
port 598 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_o[8]
port 599 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_o[9]
port 600 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 wbs_sel_i[0]
port 601 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_sel_i[1]
port 602 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 wbs_sel_i[2]
port 603 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_sel_i[3]
port 604 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_stb_i
port 605 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_we_i
port 606 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 312023 314167
string LEFview TRUE
string GDS_FILE /project/openlane/accelerator_top/runs/accelerator_top/results/magic/accelerator_top.gds
string GDS_END 160518356
string GDS_START 1411156
<< end >>

