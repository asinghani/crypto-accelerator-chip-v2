magic
tech sky130A
magscale 1 2
timestamp 1636579087
<< obsli1 >>
rect 1104 1445 248952 249713
<< obsm1 >>
rect 658 1232 249214 249744
<< metal2 >>
rect 1030 251404 1086 252204
rect 3146 251404 3202 252204
rect 5354 251404 5410 252204
rect 7562 251404 7618 252204
rect 9770 251404 9826 252204
rect 11978 251404 12034 252204
rect 14186 251404 14242 252204
rect 16302 251404 16358 252204
rect 18510 251404 18566 252204
rect 20718 251404 20774 252204
rect 22926 251404 22982 252204
rect 25134 251404 25190 252204
rect 27342 251404 27398 252204
rect 29458 251404 29514 252204
rect 31666 251404 31722 252204
rect 33874 251404 33930 252204
rect 36082 251404 36138 252204
rect 38290 251404 38346 252204
rect 40498 251404 40554 252204
rect 42706 251404 42762 252204
rect 44822 251404 44878 252204
rect 47030 251404 47086 252204
rect 49238 251404 49294 252204
rect 51446 251404 51502 252204
rect 53654 251404 53710 252204
rect 55862 251404 55918 252204
rect 57978 251404 58034 252204
rect 60186 251404 60242 252204
rect 62394 251404 62450 252204
rect 64602 251404 64658 252204
rect 66810 251404 66866 252204
rect 69018 251404 69074 252204
rect 71134 251404 71190 252204
rect 73342 251404 73398 252204
rect 75550 251404 75606 252204
rect 77758 251404 77814 252204
rect 79966 251404 80022 252204
rect 82174 251404 82230 252204
rect 84382 251404 84438 252204
rect 86498 251404 86554 252204
rect 88706 251404 88762 252204
rect 90914 251404 90970 252204
rect 93122 251404 93178 252204
rect 95330 251404 95386 252204
rect 97538 251404 97594 252204
rect 99654 251404 99710 252204
rect 101862 251404 101918 252204
rect 104070 251404 104126 252204
rect 106278 251404 106334 252204
rect 108486 251404 108542 252204
rect 110694 251404 110750 252204
rect 112810 251404 112866 252204
rect 115018 251404 115074 252204
rect 117226 251404 117282 252204
rect 119434 251404 119490 252204
rect 121642 251404 121698 252204
rect 123850 251404 123906 252204
rect 126058 251404 126114 252204
rect 128174 251404 128230 252204
rect 130382 251404 130438 252204
rect 132590 251404 132646 252204
rect 134798 251404 134854 252204
rect 137006 251404 137062 252204
rect 139214 251404 139270 252204
rect 141330 251404 141386 252204
rect 143538 251404 143594 252204
rect 145746 251404 145802 252204
rect 147954 251404 148010 252204
rect 150162 251404 150218 252204
rect 152370 251404 152426 252204
rect 154486 251404 154542 252204
rect 156694 251404 156750 252204
rect 158902 251404 158958 252204
rect 161110 251404 161166 252204
rect 163318 251404 163374 252204
rect 165526 251404 165582 252204
rect 167734 251404 167790 252204
rect 169850 251404 169906 252204
rect 172058 251404 172114 252204
rect 174266 251404 174322 252204
rect 176474 251404 176530 252204
rect 178682 251404 178738 252204
rect 180890 251404 180946 252204
rect 183006 251404 183062 252204
rect 185214 251404 185270 252204
rect 187422 251404 187478 252204
rect 189630 251404 189686 252204
rect 191838 251404 191894 252204
rect 194046 251404 194102 252204
rect 196162 251404 196218 252204
rect 198370 251404 198426 252204
rect 200578 251404 200634 252204
rect 202786 251404 202842 252204
rect 204994 251404 205050 252204
rect 207202 251404 207258 252204
rect 209410 251404 209466 252204
rect 211526 251404 211582 252204
rect 213734 251404 213790 252204
rect 215942 251404 215998 252204
rect 218150 251404 218206 252204
rect 220358 251404 220414 252204
rect 222566 251404 222622 252204
rect 224682 251404 224738 252204
rect 226890 251404 226946 252204
rect 229098 251404 229154 252204
rect 231306 251404 231362 252204
rect 233514 251404 233570 252204
rect 235722 251404 235778 252204
rect 237838 251404 237894 252204
rect 240046 251404 240102 252204
rect 242254 251404 242310 252204
rect 244462 251404 244518 252204
rect 246670 251404 246726 252204
rect 248878 251404 248934 252204
rect 202 0 258 800
rect 662 0 718 800
rect 1214 0 1270 800
rect 1674 0 1730 800
rect 2226 0 2282 800
rect 2686 0 2742 800
rect 3238 0 3294 800
rect 3698 0 3754 800
rect 4250 0 4306 800
rect 4710 0 4766 800
rect 5262 0 5318 800
rect 5814 0 5870 800
rect 6274 0 6330 800
rect 6826 0 6882 800
rect 7286 0 7342 800
rect 7838 0 7894 800
rect 8298 0 8354 800
rect 8850 0 8906 800
rect 9310 0 9366 800
rect 9862 0 9918 800
rect 10322 0 10378 800
rect 10874 0 10930 800
rect 11426 0 11482 800
rect 11886 0 11942 800
rect 12438 0 12494 800
rect 12898 0 12954 800
rect 13450 0 13506 800
rect 13910 0 13966 800
rect 14462 0 14518 800
rect 14922 0 14978 800
rect 15474 0 15530 800
rect 15934 0 15990 800
rect 16486 0 16542 800
rect 17038 0 17094 800
rect 17498 0 17554 800
rect 18050 0 18106 800
rect 18510 0 18566 800
rect 19062 0 19118 800
rect 19522 0 19578 800
rect 20074 0 20130 800
rect 20534 0 20590 800
rect 21086 0 21142 800
rect 21546 0 21602 800
rect 22098 0 22154 800
rect 22650 0 22706 800
rect 23110 0 23166 800
rect 23662 0 23718 800
rect 24122 0 24178 800
rect 24674 0 24730 800
rect 25134 0 25190 800
rect 25686 0 25742 800
rect 26146 0 26202 800
rect 26698 0 26754 800
rect 27158 0 27214 800
rect 27710 0 27766 800
rect 28262 0 28318 800
rect 28722 0 28778 800
rect 29274 0 29330 800
rect 29734 0 29790 800
rect 30286 0 30342 800
rect 30746 0 30802 800
rect 31298 0 31354 800
rect 31758 0 31814 800
rect 32310 0 32366 800
rect 32862 0 32918 800
rect 33322 0 33378 800
rect 33874 0 33930 800
rect 34334 0 34390 800
rect 34886 0 34942 800
rect 35346 0 35402 800
rect 35898 0 35954 800
rect 36358 0 36414 800
rect 36910 0 36966 800
rect 37370 0 37426 800
rect 37922 0 37978 800
rect 38474 0 38530 800
rect 38934 0 38990 800
rect 39486 0 39542 800
rect 39946 0 40002 800
rect 40498 0 40554 800
rect 40958 0 41014 800
rect 41510 0 41566 800
rect 41970 0 42026 800
rect 42522 0 42578 800
rect 42982 0 43038 800
rect 43534 0 43590 800
rect 44086 0 44142 800
rect 44546 0 44602 800
rect 45098 0 45154 800
rect 45558 0 45614 800
rect 46110 0 46166 800
rect 46570 0 46626 800
rect 47122 0 47178 800
rect 47582 0 47638 800
rect 48134 0 48190 800
rect 48594 0 48650 800
rect 49146 0 49202 800
rect 49698 0 49754 800
rect 50158 0 50214 800
rect 50710 0 50766 800
rect 51170 0 51226 800
rect 51722 0 51778 800
rect 52182 0 52238 800
rect 52734 0 52790 800
rect 53194 0 53250 800
rect 53746 0 53802 800
rect 54206 0 54262 800
rect 54758 0 54814 800
rect 55310 0 55366 800
rect 55770 0 55826 800
rect 56322 0 56378 800
rect 56782 0 56838 800
rect 57334 0 57390 800
rect 57794 0 57850 800
rect 58346 0 58402 800
rect 58806 0 58862 800
rect 59358 0 59414 800
rect 59818 0 59874 800
rect 60370 0 60426 800
rect 60922 0 60978 800
rect 61382 0 61438 800
rect 61934 0 61990 800
rect 62394 0 62450 800
rect 62946 0 63002 800
rect 63406 0 63462 800
rect 63958 0 64014 800
rect 64418 0 64474 800
rect 64970 0 65026 800
rect 65522 0 65578 800
rect 65982 0 66038 800
rect 66534 0 66590 800
rect 66994 0 67050 800
rect 67546 0 67602 800
rect 68006 0 68062 800
rect 68558 0 68614 800
rect 69018 0 69074 800
rect 69570 0 69626 800
rect 70030 0 70086 800
rect 70582 0 70638 800
rect 71134 0 71190 800
rect 71594 0 71650 800
rect 72146 0 72202 800
rect 72606 0 72662 800
rect 73158 0 73214 800
rect 73618 0 73674 800
rect 74170 0 74226 800
rect 74630 0 74686 800
rect 75182 0 75238 800
rect 75642 0 75698 800
rect 76194 0 76250 800
rect 76746 0 76802 800
rect 77206 0 77262 800
rect 77758 0 77814 800
rect 78218 0 78274 800
rect 78770 0 78826 800
rect 79230 0 79286 800
rect 79782 0 79838 800
rect 80242 0 80298 800
rect 80794 0 80850 800
rect 81254 0 81310 800
rect 81806 0 81862 800
rect 82358 0 82414 800
rect 82818 0 82874 800
rect 83370 0 83426 800
rect 83830 0 83886 800
rect 84382 0 84438 800
rect 84842 0 84898 800
rect 85394 0 85450 800
rect 85854 0 85910 800
rect 86406 0 86462 800
rect 86866 0 86922 800
rect 87418 0 87474 800
rect 87970 0 88026 800
rect 88430 0 88486 800
rect 88982 0 89038 800
rect 89442 0 89498 800
rect 89994 0 90050 800
rect 90454 0 90510 800
rect 91006 0 91062 800
rect 91466 0 91522 800
rect 92018 0 92074 800
rect 92478 0 92534 800
rect 93030 0 93086 800
rect 93582 0 93638 800
rect 94042 0 94098 800
rect 94594 0 94650 800
rect 95054 0 95110 800
rect 95606 0 95662 800
rect 96066 0 96122 800
rect 96618 0 96674 800
rect 97078 0 97134 800
rect 97630 0 97686 800
rect 98182 0 98238 800
rect 98642 0 98698 800
rect 99194 0 99250 800
rect 99654 0 99710 800
rect 100206 0 100262 800
rect 100666 0 100722 800
rect 101218 0 101274 800
rect 101678 0 101734 800
rect 102230 0 102286 800
rect 102690 0 102746 800
rect 103242 0 103298 800
rect 103794 0 103850 800
rect 104254 0 104310 800
rect 104806 0 104862 800
rect 105266 0 105322 800
rect 105818 0 105874 800
rect 106278 0 106334 800
rect 106830 0 106886 800
rect 107290 0 107346 800
rect 107842 0 107898 800
rect 108302 0 108358 800
rect 108854 0 108910 800
rect 109406 0 109462 800
rect 109866 0 109922 800
rect 110418 0 110474 800
rect 110878 0 110934 800
rect 111430 0 111486 800
rect 111890 0 111946 800
rect 112442 0 112498 800
rect 112902 0 112958 800
rect 113454 0 113510 800
rect 113914 0 113970 800
rect 114466 0 114522 800
rect 115018 0 115074 800
rect 115478 0 115534 800
rect 116030 0 116086 800
rect 116490 0 116546 800
rect 117042 0 117098 800
rect 117502 0 117558 800
rect 118054 0 118110 800
rect 118514 0 118570 800
rect 119066 0 119122 800
rect 119526 0 119582 800
rect 120078 0 120134 800
rect 120630 0 120686 800
rect 121090 0 121146 800
rect 121642 0 121698 800
rect 122102 0 122158 800
rect 122654 0 122710 800
rect 123114 0 123170 800
rect 123666 0 123722 800
rect 124126 0 124182 800
rect 124678 0 124734 800
rect 125230 0 125286 800
rect 125690 0 125746 800
rect 126242 0 126298 800
rect 126702 0 126758 800
rect 127254 0 127310 800
rect 127714 0 127770 800
rect 128266 0 128322 800
rect 128726 0 128782 800
rect 129278 0 129334 800
rect 129738 0 129794 800
rect 130290 0 130346 800
rect 130842 0 130898 800
rect 131302 0 131358 800
rect 131854 0 131910 800
rect 132314 0 132370 800
rect 132866 0 132922 800
rect 133326 0 133382 800
rect 133878 0 133934 800
rect 134338 0 134394 800
rect 134890 0 134946 800
rect 135350 0 135406 800
rect 135902 0 135958 800
rect 136454 0 136510 800
rect 136914 0 136970 800
rect 137466 0 137522 800
rect 137926 0 137982 800
rect 138478 0 138534 800
rect 138938 0 138994 800
rect 139490 0 139546 800
rect 139950 0 140006 800
rect 140502 0 140558 800
rect 140962 0 141018 800
rect 141514 0 141570 800
rect 142066 0 142122 800
rect 142526 0 142582 800
rect 143078 0 143134 800
rect 143538 0 143594 800
rect 144090 0 144146 800
rect 144550 0 144606 800
rect 145102 0 145158 800
rect 145562 0 145618 800
rect 146114 0 146170 800
rect 146574 0 146630 800
rect 147126 0 147182 800
rect 147678 0 147734 800
rect 148138 0 148194 800
rect 148690 0 148746 800
rect 149150 0 149206 800
rect 149702 0 149758 800
rect 150162 0 150218 800
rect 150714 0 150770 800
rect 151174 0 151230 800
rect 151726 0 151782 800
rect 152186 0 152242 800
rect 152738 0 152794 800
rect 153290 0 153346 800
rect 153750 0 153806 800
rect 154302 0 154358 800
rect 154762 0 154818 800
rect 155314 0 155370 800
rect 155774 0 155830 800
rect 156326 0 156382 800
rect 156786 0 156842 800
rect 157338 0 157394 800
rect 157890 0 157946 800
rect 158350 0 158406 800
rect 158902 0 158958 800
rect 159362 0 159418 800
rect 159914 0 159970 800
rect 160374 0 160430 800
rect 160926 0 160982 800
rect 161386 0 161442 800
rect 161938 0 161994 800
rect 162398 0 162454 800
rect 162950 0 163006 800
rect 163502 0 163558 800
rect 163962 0 164018 800
rect 164514 0 164570 800
rect 164974 0 165030 800
rect 165526 0 165582 800
rect 165986 0 166042 800
rect 166538 0 166594 800
rect 166998 0 167054 800
rect 167550 0 167606 800
rect 168010 0 168066 800
rect 168562 0 168618 800
rect 169114 0 169170 800
rect 169574 0 169630 800
rect 170126 0 170182 800
rect 170586 0 170642 800
rect 171138 0 171194 800
rect 171598 0 171654 800
rect 172150 0 172206 800
rect 172610 0 172666 800
rect 173162 0 173218 800
rect 173622 0 173678 800
rect 174174 0 174230 800
rect 174726 0 174782 800
rect 175186 0 175242 800
rect 175738 0 175794 800
rect 176198 0 176254 800
rect 176750 0 176806 800
rect 177210 0 177266 800
rect 177762 0 177818 800
rect 178222 0 178278 800
rect 178774 0 178830 800
rect 179234 0 179290 800
rect 179786 0 179842 800
rect 180338 0 180394 800
rect 180798 0 180854 800
rect 181350 0 181406 800
rect 181810 0 181866 800
rect 182362 0 182418 800
rect 182822 0 182878 800
rect 183374 0 183430 800
rect 183834 0 183890 800
rect 184386 0 184442 800
rect 184846 0 184902 800
rect 185398 0 185454 800
rect 185950 0 186006 800
rect 186410 0 186466 800
rect 186962 0 187018 800
rect 187422 0 187478 800
rect 187974 0 188030 800
rect 188434 0 188490 800
rect 188986 0 189042 800
rect 189446 0 189502 800
rect 189998 0 190054 800
rect 190550 0 190606 800
rect 191010 0 191066 800
rect 191562 0 191618 800
rect 192022 0 192078 800
rect 192574 0 192630 800
rect 193034 0 193090 800
rect 193586 0 193642 800
rect 194046 0 194102 800
rect 194598 0 194654 800
rect 195058 0 195114 800
rect 195610 0 195666 800
rect 196162 0 196218 800
rect 196622 0 196678 800
rect 197174 0 197230 800
rect 197634 0 197690 800
rect 198186 0 198242 800
rect 198646 0 198702 800
rect 199198 0 199254 800
rect 199658 0 199714 800
rect 200210 0 200266 800
rect 200670 0 200726 800
rect 201222 0 201278 800
rect 201774 0 201830 800
rect 202234 0 202290 800
rect 202786 0 202842 800
rect 203246 0 203302 800
rect 203798 0 203854 800
rect 204258 0 204314 800
rect 204810 0 204866 800
rect 205270 0 205326 800
rect 205822 0 205878 800
rect 206282 0 206338 800
rect 206834 0 206890 800
rect 207386 0 207442 800
rect 207846 0 207902 800
rect 208398 0 208454 800
rect 208858 0 208914 800
rect 209410 0 209466 800
rect 209870 0 209926 800
rect 210422 0 210478 800
rect 210882 0 210938 800
rect 211434 0 211490 800
rect 211894 0 211950 800
rect 212446 0 212502 800
rect 212998 0 213054 800
rect 213458 0 213514 800
rect 214010 0 214066 800
rect 214470 0 214526 800
rect 215022 0 215078 800
rect 215482 0 215538 800
rect 216034 0 216090 800
rect 216494 0 216550 800
rect 217046 0 217102 800
rect 217506 0 217562 800
rect 218058 0 218114 800
rect 218610 0 218666 800
rect 219070 0 219126 800
rect 219622 0 219678 800
rect 220082 0 220138 800
rect 220634 0 220690 800
rect 221094 0 221150 800
rect 221646 0 221702 800
rect 222106 0 222162 800
rect 222658 0 222714 800
rect 223210 0 223266 800
rect 223670 0 223726 800
rect 224222 0 224278 800
rect 224682 0 224738 800
rect 225234 0 225290 800
rect 225694 0 225750 800
rect 226246 0 226302 800
rect 226706 0 226762 800
rect 227258 0 227314 800
rect 227718 0 227774 800
rect 228270 0 228326 800
rect 228822 0 228878 800
rect 229282 0 229338 800
rect 229834 0 229890 800
rect 230294 0 230350 800
rect 230846 0 230902 800
rect 231306 0 231362 800
rect 231858 0 231914 800
rect 232318 0 232374 800
rect 232870 0 232926 800
rect 233330 0 233386 800
rect 233882 0 233938 800
rect 234434 0 234490 800
rect 234894 0 234950 800
rect 235446 0 235502 800
rect 235906 0 235962 800
rect 236458 0 236514 800
rect 236918 0 236974 800
rect 237470 0 237526 800
rect 237930 0 237986 800
rect 238482 0 238538 800
rect 238942 0 238998 800
rect 239494 0 239550 800
rect 240046 0 240102 800
rect 240506 0 240562 800
rect 241058 0 241114 800
rect 241518 0 241574 800
rect 242070 0 242126 800
rect 242530 0 242586 800
rect 243082 0 243138 800
rect 243542 0 243598 800
rect 244094 0 244150 800
rect 244554 0 244610 800
rect 245106 0 245162 800
rect 245658 0 245714 800
rect 246118 0 246174 800
rect 246670 0 246726 800
rect 247130 0 247186 800
rect 247682 0 247738 800
rect 248142 0 248198 800
rect 248694 0 248750 800
rect 249154 0 249210 800
rect 249706 0 249762 800
<< obsm2 >>
rect 18 251348 974 251546
rect 1142 251348 3090 251546
rect 3258 251348 5298 251546
rect 5466 251348 7506 251546
rect 7674 251348 9714 251546
rect 9882 251348 11922 251546
rect 12090 251348 14130 251546
rect 14298 251348 16246 251546
rect 16414 251348 18454 251546
rect 18622 251348 20662 251546
rect 20830 251348 22870 251546
rect 23038 251348 25078 251546
rect 25246 251348 27286 251546
rect 27454 251348 29402 251546
rect 29570 251348 31610 251546
rect 31778 251348 33818 251546
rect 33986 251348 36026 251546
rect 36194 251348 38234 251546
rect 38402 251348 40442 251546
rect 40610 251348 42650 251546
rect 42818 251348 44766 251546
rect 44934 251348 46974 251546
rect 47142 251348 49182 251546
rect 49350 251348 51390 251546
rect 51558 251348 53598 251546
rect 53766 251348 55806 251546
rect 55974 251348 57922 251546
rect 58090 251348 60130 251546
rect 60298 251348 62338 251546
rect 62506 251348 64546 251546
rect 64714 251348 66754 251546
rect 66922 251348 68962 251546
rect 69130 251348 71078 251546
rect 71246 251348 73286 251546
rect 73454 251348 75494 251546
rect 75662 251348 77702 251546
rect 77870 251348 79910 251546
rect 80078 251348 82118 251546
rect 82286 251348 84326 251546
rect 84494 251348 86442 251546
rect 86610 251348 88650 251546
rect 88818 251348 90858 251546
rect 91026 251348 93066 251546
rect 93234 251348 95274 251546
rect 95442 251348 97482 251546
rect 97650 251348 99598 251546
rect 99766 251348 101806 251546
rect 101974 251348 104014 251546
rect 104182 251348 106222 251546
rect 106390 251348 108430 251546
rect 108598 251348 110638 251546
rect 110806 251348 112754 251546
rect 112922 251348 114962 251546
rect 115130 251348 117170 251546
rect 117338 251348 119378 251546
rect 119546 251348 121586 251546
rect 121754 251348 123794 251546
rect 123962 251348 126002 251546
rect 126170 251348 128118 251546
rect 128286 251348 130326 251546
rect 130494 251348 132534 251546
rect 132702 251348 134742 251546
rect 134910 251348 136950 251546
rect 137118 251348 139158 251546
rect 139326 251348 141274 251546
rect 141442 251348 143482 251546
rect 143650 251348 145690 251546
rect 145858 251348 147898 251546
rect 148066 251348 150106 251546
rect 150274 251348 152314 251546
rect 152482 251348 154430 251546
rect 154598 251348 156638 251546
rect 156806 251348 158846 251546
rect 159014 251348 161054 251546
rect 161222 251348 163262 251546
rect 163430 251348 165470 251546
rect 165638 251348 167678 251546
rect 167846 251348 169794 251546
rect 169962 251348 172002 251546
rect 172170 251348 174210 251546
rect 174378 251348 176418 251546
rect 176586 251348 178626 251546
rect 178794 251348 180834 251546
rect 181002 251348 182950 251546
rect 183118 251348 185158 251546
rect 185326 251348 187366 251546
rect 187534 251348 189574 251546
rect 189742 251348 191782 251546
rect 191950 251348 193990 251546
rect 194158 251348 196106 251546
rect 196274 251348 198314 251546
rect 198482 251348 200522 251546
rect 200690 251348 202730 251546
rect 202898 251348 204938 251546
rect 205106 251348 207146 251546
rect 207314 251348 209354 251546
rect 209522 251348 211470 251546
rect 211638 251348 213678 251546
rect 213846 251348 215886 251546
rect 216054 251348 218094 251546
rect 218262 251348 220302 251546
rect 220470 251348 222510 251546
rect 222678 251348 224626 251546
rect 224794 251348 226834 251546
rect 227002 251348 229042 251546
rect 229210 251348 231250 251546
rect 231418 251348 233458 251546
rect 233626 251348 235666 251546
rect 235834 251348 237782 251546
rect 237950 251348 239990 251546
rect 240158 251348 242198 251546
rect 242366 251348 244406 251546
rect 244574 251348 246614 251546
rect 246782 251348 248822 251546
rect 248990 251348 249208 251546
rect 18 856 249208 251348
rect 18 734 146 856
rect 314 734 606 856
rect 774 734 1158 856
rect 1326 734 1618 856
rect 1786 734 2170 856
rect 2338 734 2630 856
rect 2798 734 3182 856
rect 3350 734 3642 856
rect 3810 734 4194 856
rect 4362 734 4654 856
rect 4822 734 5206 856
rect 5374 734 5758 856
rect 5926 734 6218 856
rect 6386 734 6770 856
rect 6938 734 7230 856
rect 7398 734 7782 856
rect 7950 734 8242 856
rect 8410 734 8794 856
rect 8962 734 9254 856
rect 9422 734 9806 856
rect 9974 734 10266 856
rect 10434 734 10818 856
rect 10986 734 11370 856
rect 11538 734 11830 856
rect 11998 734 12382 856
rect 12550 734 12842 856
rect 13010 734 13394 856
rect 13562 734 13854 856
rect 14022 734 14406 856
rect 14574 734 14866 856
rect 15034 734 15418 856
rect 15586 734 15878 856
rect 16046 734 16430 856
rect 16598 734 16982 856
rect 17150 734 17442 856
rect 17610 734 17994 856
rect 18162 734 18454 856
rect 18622 734 19006 856
rect 19174 734 19466 856
rect 19634 734 20018 856
rect 20186 734 20478 856
rect 20646 734 21030 856
rect 21198 734 21490 856
rect 21658 734 22042 856
rect 22210 734 22594 856
rect 22762 734 23054 856
rect 23222 734 23606 856
rect 23774 734 24066 856
rect 24234 734 24618 856
rect 24786 734 25078 856
rect 25246 734 25630 856
rect 25798 734 26090 856
rect 26258 734 26642 856
rect 26810 734 27102 856
rect 27270 734 27654 856
rect 27822 734 28206 856
rect 28374 734 28666 856
rect 28834 734 29218 856
rect 29386 734 29678 856
rect 29846 734 30230 856
rect 30398 734 30690 856
rect 30858 734 31242 856
rect 31410 734 31702 856
rect 31870 734 32254 856
rect 32422 734 32806 856
rect 32974 734 33266 856
rect 33434 734 33818 856
rect 33986 734 34278 856
rect 34446 734 34830 856
rect 34998 734 35290 856
rect 35458 734 35842 856
rect 36010 734 36302 856
rect 36470 734 36854 856
rect 37022 734 37314 856
rect 37482 734 37866 856
rect 38034 734 38418 856
rect 38586 734 38878 856
rect 39046 734 39430 856
rect 39598 734 39890 856
rect 40058 734 40442 856
rect 40610 734 40902 856
rect 41070 734 41454 856
rect 41622 734 41914 856
rect 42082 734 42466 856
rect 42634 734 42926 856
rect 43094 734 43478 856
rect 43646 734 44030 856
rect 44198 734 44490 856
rect 44658 734 45042 856
rect 45210 734 45502 856
rect 45670 734 46054 856
rect 46222 734 46514 856
rect 46682 734 47066 856
rect 47234 734 47526 856
rect 47694 734 48078 856
rect 48246 734 48538 856
rect 48706 734 49090 856
rect 49258 734 49642 856
rect 49810 734 50102 856
rect 50270 734 50654 856
rect 50822 734 51114 856
rect 51282 734 51666 856
rect 51834 734 52126 856
rect 52294 734 52678 856
rect 52846 734 53138 856
rect 53306 734 53690 856
rect 53858 734 54150 856
rect 54318 734 54702 856
rect 54870 734 55254 856
rect 55422 734 55714 856
rect 55882 734 56266 856
rect 56434 734 56726 856
rect 56894 734 57278 856
rect 57446 734 57738 856
rect 57906 734 58290 856
rect 58458 734 58750 856
rect 58918 734 59302 856
rect 59470 734 59762 856
rect 59930 734 60314 856
rect 60482 734 60866 856
rect 61034 734 61326 856
rect 61494 734 61878 856
rect 62046 734 62338 856
rect 62506 734 62890 856
rect 63058 734 63350 856
rect 63518 734 63902 856
rect 64070 734 64362 856
rect 64530 734 64914 856
rect 65082 734 65466 856
rect 65634 734 65926 856
rect 66094 734 66478 856
rect 66646 734 66938 856
rect 67106 734 67490 856
rect 67658 734 67950 856
rect 68118 734 68502 856
rect 68670 734 68962 856
rect 69130 734 69514 856
rect 69682 734 69974 856
rect 70142 734 70526 856
rect 70694 734 71078 856
rect 71246 734 71538 856
rect 71706 734 72090 856
rect 72258 734 72550 856
rect 72718 734 73102 856
rect 73270 734 73562 856
rect 73730 734 74114 856
rect 74282 734 74574 856
rect 74742 734 75126 856
rect 75294 734 75586 856
rect 75754 734 76138 856
rect 76306 734 76690 856
rect 76858 734 77150 856
rect 77318 734 77702 856
rect 77870 734 78162 856
rect 78330 734 78714 856
rect 78882 734 79174 856
rect 79342 734 79726 856
rect 79894 734 80186 856
rect 80354 734 80738 856
rect 80906 734 81198 856
rect 81366 734 81750 856
rect 81918 734 82302 856
rect 82470 734 82762 856
rect 82930 734 83314 856
rect 83482 734 83774 856
rect 83942 734 84326 856
rect 84494 734 84786 856
rect 84954 734 85338 856
rect 85506 734 85798 856
rect 85966 734 86350 856
rect 86518 734 86810 856
rect 86978 734 87362 856
rect 87530 734 87914 856
rect 88082 734 88374 856
rect 88542 734 88926 856
rect 89094 734 89386 856
rect 89554 734 89938 856
rect 90106 734 90398 856
rect 90566 734 90950 856
rect 91118 734 91410 856
rect 91578 734 91962 856
rect 92130 734 92422 856
rect 92590 734 92974 856
rect 93142 734 93526 856
rect 93694 734 93986 856
rect 94154 734 94538 856
rect 94706 734 94998 856
rect 95166 734 95550 856
rect 95718 734 96010 856
rect 96178 734 96562 856
rect 96730 734 97022 856
rect 97190 734 97574 856
rect 97742 734 98126 856
rect 98294 734 98586 856
rect 98754 734 99138 856
rect 99306 734 99598 856
rect 99766 734 100150 856
rect 100318 734 100610 856
rect 100778 734 101162 856
rect 101330 734 101622 856
rect 101790 734 102174 856
rect 102342 734 102634 856
rect 102802 734 103186 856
rect 103354 734 103738 856
rect 103906 734 104198 856
rect 104366 734 104750 856
rect 104918 734 105210 856
rect 105378 734 105762 856
rect 105930 734 106222 856
rect 106390 734 106774 856
rect 106942 734 107234 856
rect 107402 734 107786 856
rect 107954 734 108246 856
rect 108414 734 108798 856
rect 108966 734 109350 856
rect 109518 734 109810 856
rect 109978 734 110362 856
rect 110530 734 110822 856
rect 110990 734 111374 856
rect 111542 734 111834 856
rect 112002 734 112386 856
rect 112554 734 112846 856
rect 113014 734 113398 856
rect 113566 734 113858 856
rect 114026 734 114410 856
rect 114578 734 114962 856
rect 115130 734 115422 856
rect 115590 734 115974 856
rect 116142 734 116434 856
rect 116602 734 116986 856
rect 117154 734 117446 856
rect 117614 734 117998 856
rect 118166 734 118458 856
rect 118626 734 119010 856
rect 119178 734 119470 856
rect 119638 734 120022 856
rect 120190 734 120574 856
rect 120742 734 121034 856
rect 121202 734 121586 856
rect 121754 734 122046 856
rect 122214 734 122598 856
rect 122766 734 123058 856
rect 123226 734 123610 856
rect 123778 734 124070 856
rect 124238 734 124622 856
rect 124790 734 125174 856
rect 125342 734 125634 856
rect 125802 734 126186 856
rect 126354 734 126646 856
rect 126814 734 127198 856
rect 127366 734 127658 856
rect 127826 734 128210 856
rect 128378 734 128670 856
rect 128838 734 129222 856
rect 129390 734 129682 856
rect 129850 734 130234 856
rect 130402 734 130786 856
rect 130954 734 131246 856
rect 131414 734 131798 856
rect 131966 734 132258 856
rect 132426 734 132810 856
rect 132978 734 133270 856
rect 133438 734 133822 856
rect 133990 734 134282 856
rect 134450 734 134834 856
rect 135002 734 135294 856
rect 135462 734 135846 856
rect 136014 734 136398 856
rect 136566 734 136858 856
rect 137026 734 137410 856
rect 137578 734 137870 856
rect 138038 734 138422 856
rect 138590 734 138882 856
rect 139050 734 139434 856
rect 139602 734 139894 856
rect 140062 734 140446 856
rect 140614 734 140906 856
rect 141074 734 141458 856
rect 141626 734 142010 856
rect 142178 734 142470 856
rect 142638 734 143022 856
rect 143190 734 143482 856
rect 143650 734 144034 856
rect 144202 734 144494 856
rect 144662 734 145046 856
rect 145214 734 145506 856
rect 145674 734 146058 856
rect 146226 734 146518 856
rect 146686 734 147070 856
rect 147238 734 147622 856
rect 147790 734 148082 856
rect 148250 734 148634 856
rect 148802 734 149094 856
rect 149262 734 149646 856
rect 149814 734 150106 856
rect 150274 734 150658 856
rect 150826 734 151118 856
rect 151286 734 151670 856
rect 151838 734 152130 856
rect 152298 734 152682 856
rect 152850 734 153234 856
rect 153402 734 153694 856
rect 153862 734 154246 856
rect 154414 734 154706 856
rect 154874 734 155258 856
rect 155426 734 155718 856
rect 155886 734 156270 856
rect 156438 734 156730 856
rect 156898 734 157282 856
rect 157450 734 157834 856
rect 158002 734 158294 856
rect 158462 734 158846 856
rect 159014 734 159306 856
rect 159474 734 159858 856
rect 160026 734 160318 856
rect 160486 734 160870 856
rect 161038 734 161330 856
rect 161498 734 161882 856
rect 162050 734 162342 856
rect 162510 734 162894 856
rect 163062 734 163446 856
rect 163614 734 163906 856
rect 164074 734 164458 856
rect 164626 734 164918 856
rect 165086 734 165470 856
rect 165638 734 165930 856
rect 166098 734 166482 856
rect 166650 734 166942 856
rect 167110 734 167494 856
rect 167662 734 167954 856
rect 168122 734 168506 856
rect 168674 734 169058 856
rect 169226 734 169518 856
rect 169686 734 170070 856
rect 170238 734 170530 856
rect 170698 734 171082 856
rect 171250 734 171542 856
rect 171710 734 172094 856
rect 172262 734 172554 856
rect 172722 734 173106 856
rect 173274 734 173566 856
rect 173734 734 174118 856
rect 174286 734 174670 856
rect 174838 734 175130 856
rect 175298 734 175682 856
rect 175850 734 176142 856
rect 176310 734 176694 856
rect 176862 734 177154 856
rect 177322 734 177706 856
rect 177874 734 178166 856
rect 178334 734 178718 856
rect 178886 734 179178 856
rect 179346 734 179730 856
rect 179898 734 180282 856
rect 180450 734 180742 856
rect 180910 734 181294 856
rect 181462 734 181754 856
rect 181922 734 182306 856
rect 182474 734 182766 856
rect 182934 734 183318 856
rect 183486 734 183778 856
rect 183946 734 184330 856
rect 184498 734 184790 856
rect 184958 734 185342 856
rect 185510 734 185894 856
rect 186062 734 186354 856
rect 186522 734 186906 856
rect 187074 734 187366 856
rect 187534 734 187918 856
rect 188086 734 188378 856
rect 188546 734 188930 856
rect 189098 734 189390 856
rect 189558 734 189942 856
rect 190110 734 190494 856
rect 190662 734 190954 856
rect 191122 734 191506 856
rect 191674 734 191966 856
rect 192134 734 192518 856
rect 192686 734 192978 856
rect 193146 734 193530 856
rect 193698 734 193990 856
rect 194158 734 194542 856
rect 194710 734 195002 856
rect 195170 734 195554 856
rect 195722 734 196106 856
rect 196274 734 196566 856
rect 196734 734 197118 856
rect 197286 734 197578 856
rect 197746 734 198130 856
rect 198298 734 198590 856
rect 198758 734 199142 856
rect 199310 734 199602 856
rect 199770 734 200154 856
rect 200322 734 200614 856
rect 200782 734 201166 856
rect 201334 734 201718 856
rect 201886 734 202178 856
rect 202346 734 202730 856
rect 202898 734 203190 856
rect 203358 734 203742 856
rect 203910 734 204202 856
rect 204370 734 204754 856
rect 204922 734 205214 856
rect 205382 734 205766 856
rect 205934 734 206226 856
rect 206394 734 206778 856
rect 206946 734 207330 856
rect 207498 734 207790 856
rect 207958 734 208342 856
rect 208510 734 208802 856
rect 208970 734 209354 856
rect 209522 734 209814 856
rect 209982 734 210366 856
rect 210534 734 210826 856
rect 210994 734 211378 856
rect 211546 734 211838 856
rect 212006 734 212390 856
rect 212558 734 212942 856
rect 213110 734 213402 856
rect 213570 734 213954 856
rect 214122 734 214414 856
rect 214582 734 214966 856
rect 215134 734 215426 856
rect 215594 734 215978 856
rect 216146 734 216438 856
rect 216606 734 216990 856
rect 217158 734 217450 856
rect 217618 734 218002 856
rect 218170 734 218554 856
rect 218722 734 219014 856
rect 219182 734 219566 856
rect 219734 734 220026 856
rect 220194 734 220578 856
rect 220746 734 221038 856
rect 221206 734 221590 856
rect 221758 734 222050 856
rect 222218 734 222602 856
rect 222770 734 223154 856
rect 223322 734 223614 856
rect 223782 734 224166 856
rect 224334 734 224626 856
rect 224794 734 225178 856
rect 225346 734 225638 856
rect 225806 734 226190 856
rect 226358 734 226650 856
rect 226818 734 227202 856
rect 227370 734 227662 856
rect 227830 734 228214 856
rect 228382 734 228766 856
rect 228934 734 229226 856
rect 229394 734 229778 856
rect 229946 734 230238 856
rect 230406 734 230790 856
rect 230958 734 231250 856
rect 231418 734 231802 856
rect 231970 734 232262 856
rect 232430 734 232814 856
rect 232982 734 233274 856
rect 233442 734 233826 856
rect 233994 734 234378 856
rect 234546 734 234838 856
rect 235006 734 235390 856
rect 235558 734 235850 856
rect 236018 734 236402 856
rect 236570 734 236862 856
rect 237030 734 237414 856
rect 237582 734 237874 856
rect 238042 734 238426 856
rect 238594 734 238886 856
rect 239054 734 239438 856
rect 239606 734 239990 856
rect 240158 734 240450 856
rect 240618 734 241002 856
rect 241170 734 241462 856
rect 241630 734 242014 856
rect 242182 734 242474 856
rect 242642 734 243026 856
rect 243194 734 243486 856
rect 243654 734 244038 856
rect 244206 734 244498 856
rect 244666 734 245050 856
rect 245218 734 245602 856
rect 245770 734 246062 856
rect 246230 734 246614 856
rect 246782 734 247074 856
rect 247242 734 247626 856
rect 247794 734 248086 856
rect 248254 734 248638 856
rect 248806 734 249098 856
<< obsm3 >>
rect 13 1939 246087 249729
<< metal4 >>
rect 4208 2128 4528 249744
rect 19568 2128 19888 249744
rect 34928 2128 35248 249744
rect 50288 2128 50608 249744
rect 65648 2128 65968 249744
rect 81008 2128 81328 249744
rect 96368 2128 96688 249744
rect 111728 2128 112048 249744
rect 127088 2128 127408 249744
rect 142448 2128 142768 249744
rect 157808 2128 158128 249744
rect 173168 2128 173488 249744
rect 188528 2128 188848 249744
rect 203888 2128 204208 249744
rect 219248 2128 219568 249744
rect 234608 2128 234928 249744
<< obsm4 >>
rect 16803 3027 19488 248437
rect 19968 3027 34848 248437
rect 35328 3027 50208 248437
rect 50688 3027 65568 248437
rect 66048 3027 80928 248437
rect 81408 3027 96288 248437
rect 96768 3027 111648 248437
rect 112128 3027 127008 248437
rect 127488 3027 142368 248437
rect 142848 3027 157728 248437
rect 158208 3027 173088 248437
rect 173568 3027 188448 248437
rect 188928 3027 203808 248437
rect 204288 3027 219168 248437
rect 219648 3027 234528 248437
rect 235008 3027 236749 248437
<< labels >>
rlabel metal2 s 1030 251404 1086 252204 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 66810 251404 66866 252204 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 73342 251404 73398 252204 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 79966 251404 80022 252204 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 86498 251404 86554 252204 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 93122 251404 93178 252204 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 99654 251404 99710 252204 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 106278 251404 106334 252204 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 112810 251404 112866 252204 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 119434 251404 119490 252204 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 126058 251404 126114 252204 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 7562 251404 7618 252204 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 132590 251404 132646 252204 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 139214 251404 139270 252204 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 145746 251404 145802 252204 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 152370 251404 152426 252204 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 158902 251404 158958 252204 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 165526 251404 165582 252204 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 172058 251404 172114 252204 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 178682 251404 178738 252204 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 185214 251404 185270 252204 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 191838 251404 191894 252204 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 14186 251404 14242 252204 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 198370 251404 198426 252204 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 204994 251404 205050 252204 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 211526 251404 211582 252204 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 218150 251404 218206 252204 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 224682 251404 224738 252204 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 231306 251404 231362 252204 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 237838 251404 237894 252204 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 244462 251404 244518 252204 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 20718 251404 20774 252204 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 27342 251404 27398 252204 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 33874 251404 33930 252204 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 40498 251404 40554 252204 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 47030 251404 47086 252204 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 53654 251404 53710 252204 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 60186 251404 60242 252204 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3146 251404 3202 252204 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 69018 251404 69074 252204 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 75550 251404 75606 252204 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 82174 251404 82230 252204 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 88706 251404 88762 252204 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 95330 251404 95386 252204 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 101862 251404 101918 252204 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 108486 251404 108542 252204 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 115018 251404 115074 252204 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 121642 251404 121698 252204 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 128174 251404 128230 252204 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 9770 251404 9826 252204 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 134798 251404 134854 252204 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 141330 251404 141386 252204 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 147954 251404 148010 252204 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 154486 251404 154542 252204 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 161110 251404 161166 252204 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 167734 251404 167790 252204 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 174266 251404 174322 252204 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 180890 251404 180946 252204 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 187422 251404 187478 252204 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 194046 251404 194102 252204 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 16302 251404 16358 252204 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 200578 251404 200634 252204 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 207202 251404 207258 252204 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 213734 251404 213790 252204 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 220358 251404 220414 252204 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 226890 251404 226946 252204 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 233514 251404 233570 252204 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 240046 251404 240102 252204 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 246670 251404 246726 252204 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 22926 251404 22982 252204 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 29458 251404 29514 252204 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 36082 251404 36138 252204 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 42706 251404 42762 252204 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 49238 251404 49294 252204 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 55862 251404 55918 252204 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 62394 251404 62450 252204 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 5354 251404 5410 252204 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 71134 251404 71190 252204 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 77758 251404 77814 252204 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 84382 251404 84438 252204 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 90914 251404 90970 252204 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 97538 251404 97594 252204 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 104070 251404 104126 252204 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 110694 251404 110750 252204 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 117226 251404 117282 252204 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 123850 251404 123906 252204 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 130382 251404 130438 252204 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 11978 251404 12034 252204 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 137006 251404 137062 252204 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 143538 251404 143594 252204 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 150162 251404 150218 252204 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 156694 251404 156750 252204 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 163318 251404 163374 252204 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 169850 251404 169906 252204 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 176474 251404 176530 252204 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 183006 251404 183062 252204 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 189630 251404 189686 252204 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 196162 251404 196218 252204 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 18510 251404 18566 252204 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 202786 251404 202842 252204 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 209410 251404 209466 252204 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 215942 251404 215998 252204 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 222566 251404 222622 252204 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 229098 251404 229154 252204 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 235722 251404 235778 252204 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 242254 251404 242310 252204 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 248878 251404 248934 252204 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 25134 251404 25190 252204 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 31666 251404 31722 252204 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 38290 251404 38346 252204 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 44822 251404 44878 252204 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 51446 251404 51502 252204 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 57978 251404 58034 252204 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 64602 251404 64658 252204 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 54206 0 54262 800 6 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 207386 0 207442 800 6 la_data_in[100]
port 116 nsew signal input
rlabel metal2 s 208858 0 208914 800 6 la_data_in[101]
port 117 nsew signal input
rlabel metal2 s 210422 0 210478 800 6 la_data_in[102]
port 118 nsew signal input
rlabel metal2 s 211894 0 211950 800 6 la_data_in[103]
port 119 nsew signal input
rlabel metal2 s 213458 0 213514 800 6 la_data_in[104]
port 120 nsew signal input
rlabel metal2 s 215022 0 215078 800 6 la_data_in[105]
port 121 nsew signal input
rlabel metal2 s 216494 0 216550 800 6 la_data_in[106]
port 122 nsew signal input
rlabel metal2 s 218058 0 218114 800 6 la_data_in[107]
port 123 nsew signal input
rlabel metal2 s 219622 0 219678 800 6 la_data_in[108]
port 124 nsew signal input
rlabel metal2 s 221094 0 221150 800 6 la_data_in[109]
port 125 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_data_in[10]
port 126 nsew signal input
rlabel metal2 s 222658 0 222714 800 6 la_data_in[110]
port 127 nsew signal input
rlabel metal2 s 224222 0 224278 800 6 la_data_in[111]
port 128 nsew signal input
rlabel metal2 s 225694 0 225750 800 6 la_data_in[112]
port 129 nsew signal input
rlabel metal2 s 227258 0 227314 800 6 la_data_in[113]
port 130 nsew signal input
rlabel metal2 s 228822 0 228878 800 6 la_data_in[114]
port 131 nsew signal input
rlabel metal2 s 230294 0 230350 800 6 la_data_in[115]
port 132 nsew signal input
rlabel metal2 s 231858 0 231914 800 6 la_data_in[116]
port 133 nsew signal input
rlabel metal2 s 233330 0 233386 800 6 la_data_in[117]
port 134 nsew signal input
rlabel metal2 s 234894 0 234950 800 6 la_data_in[118]
port 135 nsew signal input
rlabel metal2 s 236458 0 236514 800 6 la_data_in[119]
port 136 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_data_in[11]
port 137 nsew signal input
rlabel metal2 s 237930 0 237986 800 6 la_data_in[120]
port 138 nsew signal input
rlabel metal2 s 239494 0 239550 800 6 la_data_in[121]
port 139 nsew signal input
rlabel metal2 s 241058 0 241114 800 6 la_data_in[122]
port 140 nsew signal input
rlabel metal2 s 242530 0 242586 800 6 la_data_in[123]
port 141 nsew signal input
rlabel metal2 s 244094 0 244150 800 6 la_data_in[124]
port 142 nsew signal input
rlabel metal2 s 245658 0 245714 800 6 la_data_in[125]
port 143 nsew signal input
rlabel metal2 s 247130 0 247186 800 6 la_data_in[126]
port 144 nsew signal input
rlabel metal2 s 248694 0 248750 800 6 la_data_in[127]
port 145 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 la_data_in[12]
port 146 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 la_data_in[13]
port 147 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 la_data_in[14]
port 148 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_data_in[15]
port 149 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_data_in[16]
port 150 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 la_data_in[17]
port 151 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_data_in[18]
port 152 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 la_data_in[19]
port 153 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 la_data_in[1]
port 154 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_data_in[20]
port 155 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 la_data_in[21]
port 156 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_data_in[22]
port 157 nsew signal input
rlabel metal2 s 89442 0 89498 800 6 la_data_in[23]
port 158 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 la_data_in[24]
port 159 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 la_data_in[25]
port 160 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_data_in[26]
port 161 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 la_data_in[27]
port 162 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_data_in[28]
port 163 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_data_in[29]
port 164 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_data_in[2]
port 165 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 la_data_in[30]
port 166 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_data_in[31]
port 167 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_data_in[32]
port 168 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_data_in[33]
port 169 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 la_data_in[34]
port 170 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 la_data_in[35]
port 171 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 la_data_in[36]
port 172 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 la_data_in[37]
port 173 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_data_in[38]
port 174 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 la_data_in[39]
port 175 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_data_in[3]
port 176 nsew signal input
rlabel metal2 s 115478 0 115534 800 6 la_data_in[40]
port 177 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 la_data_in[41]
port 178 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 la_data_in[42]
port 179 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 la_data_in[43]
port 180 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 la_data_in[44]
port 181 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 la_data_in[45]
port 182 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 la_data_in[46]
port 183 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 la_data_in[47]
port 184 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 la_data_in[48]
port 185 nsew signal input
rlabel metal2 s 129278 0 129334 800 6 la_data_in[49]
port 186 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 la_data_in[4]
port 187 nsew signal input
rlabel metal2 s 130842 0 130898 800 6 la_data_in[50]
port 188 nsew signal input
rlabel metal2 s 132314 0 132370 800 6 la_data_in[51]
port 189 nsew signal input
rlabel metal2 s 133878 0 133934 800 6 la_data_in[52]
port 190 nsew signal input
rlabel metal2 s 135350 0 135406 800 6 la_data_in[53]
port 191 nsew signal input
rlabel metal2 s 136914 0 136970 800 6 la_data_in[54]
port 192 nsew signal input
rlabel metal2 s 138478 0 138534 800 6 la_data_in[55]
port 193 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 la_data_in[56]
port 194 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 la_data_in[57]
port 195 nsew signal input
rlabel metal2 s 143078 0 143134 800 6 la_data_in[58]
port 196 nsew signal input
rlabel metal2 s 144550 0 144606 800 6 la_data_in[59]
port 197 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 la_data_in[5]
port 198 nsew signal input
rlabel metal2 s 146114 0 146170 800 6 la_data_in[60]
port 199 nsew signal input
rlabel metal2 s 147678 0 147734 800 6 la_data_in[61]
port 200 nsew signal input
rlabel metal2 s 149150 0 149206 800 6 la_data_in[62]
port 201 nsew signal input
rlabel metal2 s 150714 0 150770 800 6 la_data_in[63]
port 202 nsew signal input
rlabel metal2 s 152186 0 152242 800 6 la_data_in[64]
port 203 nsew signal input
rlabel metal2 s 153750 0 153806 800 6 la_data_in[65]
port 204 nsew signal input
rlabel metal2 s 155314 0 155370 800 6 la_data_in[66]
port 205 nsew signal input
rlabel metal2 s 156786 0 156842 800 6 la_data_in[67]
port 206 nsew signal input
rlabel metal2 s 158350 0 158406 800 6 la_data_in[68]
port 207 nsew signal input
rlabel metal2 s 159914 0 159970 800 6 la_data_in[69]
port 208 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_data_in[6]
port 209 nsew signal input
rlabel metal2 s 161386 0 161442 800 6 la_data_in[70]
port 210 nsew signal input
rlabel metal2 s 162950 0 163006 800 6 la_data_in[71]
port 211 nsew signal input
rlabel metal2 s 164514 0 164570 800 6 la_data_in[72]
port 212 nsew signal input
rlabel metal2 s 165986 0 166042 800 6 la_data_in[73]
port 213 nsew signal input
rlabel metal2 s 167550 0 167606 800 6 la_data_in[74]
port 214 nsew signal input
rlabel metal2 s 169114 0 169170 800 6 la_data_in[75]
port 215 nsew signal input
rlabel metal2 s 170586 0 170642 800 6 la_data_in[76]
port 216 nsew signal input
rlabel metal2 s 172150 0 172206 800 6 la_data_in[77]
port 217 nsew signal input
rlabel metal2 s 173622 0 173678 800 6 la_data_in[78]
port 218 nsew signal input
rlabel metal2 s 175186 0 175242 800 6 la_data_in[79]
port 219 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 la_data_in[7]
port 220 nsew signal input
rlabel metal2 s 176750 0 176806 800 6 la_data_in[80]
port 221 nsew signal input
rlabel metal2 s 178222 0 178278 800 6 la_data_in[81]
port 222 nsew signal input
rlabel metal2 s 179786 0 179842 800 6 la_data_in[82]
port 223 nsew signal input
rlabel metal2 s 181350 0 181406 800 6 la_data_in[83]
port 224 nsew signal input
rlabel metal2 s 182822 0 182878 800 6 la_data_in[84]
port 225 nsew signal input
rlabel metal2 s 184386 0 184442 800 6 la_data_in[85]
port 226 nsew signal input
rlabel metal2 s 185950 0 186006 800 6 la_data_in[86]
port 227 nsew signal input
rlabel metal2 s 187422 0 187478 800 6 la_data_in[87]
port 228 nsew signal input
rlabel metal2 s 188986 0 189042 800 6 la_data_in[88]
port 229 nsew signal input
rlabel metal2 s 190550 0 190606 800 6 la_data_in[89]
port 230 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_data_in[8]
port 231 nsew signal input
rlabel metal2 s 192022 0 192078 800 6 la_data_in[90]
port 232 nsew signal input
rlabel metal2 s 193586 0 193642 800 6 la_data_in[91]
port 233 nsew signal input
rlabel metal2 s 195058 0 195114 800 6 la_data_in[92]
port 234 nsew signal input
rlabel metal2 s 196622 0 196678 800 6 la_data_in[93]
port 235 nsew signal input
rlabel metal2 s 198186 0 198242 800 6 la_data_in[94]
port 236 nsew signal input
rlabel metal2 s 199658 0 199714 800 6 la_data_in[95]
port 237 nsew signal input
rlabel metal2 s 201222 0 201278 800 6 la_data_in[96]
port 238 nsew signal input
rlabel metal2 s 202786 0 202842 800 6 la_data_in[97]
port 239 nsew signal input
rlabel metal2 s 204258 0 204314 800 6 la_data_in[98]
port 240 nsew signal input
rlabel metal2 s 205822 0 205878 800 6 la_data_in[99]
port 241 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 la_data_in[9]
port 242 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 la_data_out[0]
port 243 nsew signal output
rlabel metal2 s 207846 0 207902 800 6 la_data_out[100]
port 244 nsew signal output
rlabel metal2 s 209410 0 209466 800 6 la_data_out[101]
port 245 nsew signal output
rlabel metal2 s 210882 0 210938 800 6 la_data_out[102]
port 246 nsew signal output
rlabel metal2 s 212446 0 212502 800 6 la_data_out[103]
port 247 nsew signal output
rlabel metal2 s 214010 0 214066 800 6 la_data_out[104]
port 248 nsew signal output
rlabel metal2 s 215482 0 215538 800 6 la_data_out[105]
port 249 nsew signal output
rlabel metal2 s 217046 0 217102 800 6 la_data_out[106]
port 250 nsew signal output
rlabel metal2 s 218610 0 218666 800 6 la_data_out[107]
port 251 nsew signal output
rlabel metal2 s 220082 0 220138 800 6 la_data_out[108]
port 252 nsew signal output
rlabel metal2 s 221646 0 221702 800 6 la_data_out[109]
port 253 nsew signal output
rlabel metal2 s 70030 0 70086 800 6 la_data_out[10]
port 254 nsew signal output
rlabel metal2 s 223210 0 223266 800 6 la_data_out[110]
port 255 nsew signal output
rlabel metal2 s 224682 0 224738 800 6 la_data_out[111]
port 256 nsew signal output
rlabel metal2 s 226246 0 226302 800 6 la_data_out[112]
port 257 nsew signal output
rlabel metal2 s 227718 0 227774 800 6 la_data_out[113]
port 258 nsew signal output
rlabel metal2 s 229282 0 229338 800 6 la_data_out[114]
port 259 nsew signal output
rlabel metal2 s 230846 0 230902 800 6 la_data_out[115]
port 260 nsew signal output
rlabel metal2 s 232318 0 232374 800 6 la_data_out[116]
port 261 nsew signal output
rlabel metal2 s 233882 0 233938 800 6 la_data_out[117]
port 262 nsew signal output
rlabel metal2 s 235446 0 235502 800 6 la_data_out[118]
port 263 nsew signal output
rlabel metal2 s 236918 0 236974 800 6 la_data_out[119]
port 264 nsew signal output
rlabel metal2 s 71594 0 71650 800 6 la_data_out[11]
port 265 nsew signal output
rlabel metal2 s 238482 0 238538 800 6 la_data_out[120]
port 266 nsew signal output
rlabel metal2 s 240046 0 240102 800 6 la_data_out[121]
port 267 nsew signal output
rlabel metal2 s 241518 0 241574 800 6 la_data_out[122]
port 268 nsew signal output
rlabel metal2 s 243082 0 243138 800 6 la_data_out[123]
port 269 nsew signal output
rlabel metal2 s 244554 0 244610 800 6 la_data_out[124]
port 270 nsew signal output
rlabel metal2 s 246118 0 246174 800 6 la_data_out[125]
port 271 nsew signal output
rlabel metal2 s 247682 0 247738 800 6 la_data_out[126]
port 272 nsew signal output
rlabel metal2 s 249154 0 249210 800 6 la_data_out[127]
port 273 nsew signal output
rlabel metal2 s 73158 0 73214 800 6 la_data_out[12]
port 274 nsew signal output
rlabel metal2 s 74630 0 74686 800 6 la_data_out[13]
port 275 nsew signal output
rlabel metal2 s 76194 0 76250 800 6 la_data_out[14]
port 276 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 la_data_out[15]
port 277 nsew signal output
rlabel metal2 s 79230 0 79286 800 6 la_data_out[16]
port 278 nsew signal output
rlabel metal2 s 80794 0 80850 800 6 la_data_out[17]
port 279 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 la_data_out[18]
port 280 nsew signal output
rlabel metal2 s 83830 0 83886 800 6 la_data_out[19]
port 281 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 la_data_out[1]
port 282 nsew signal output
rlabel metal2 s 85394 0 85450 800 6 la_data_out[20]
port 283 nsew signal output
rlabel metal2 s 86866 0 86922 800 6 la_data_out[21]
port 284 nsew signal output
rlabel metal2 s 88430 0 88486 800 6 la_data_out[22]
port 285 nsew signal output
rlabel metal2 s 89994 0 90050 800 6 la_data_out[23]
port 286 nsew signal output
rlabel metal2 s 91466 0 91522 800 6 la_data_out[24]
port 287 nsew signal output
rlabel metal2 s 93030 0 93086 800 6 la_data_out[25]
port 288 nsew signal output
rlabel metal2 s 94594 0 94650 800 6 la_data_out[26]
port 289 nsew signal output
rlabel metal2 s 96066 0 96122 800 6 la_data_out[27]
port 290 nsew signal output
rlabel metal2 s 97630 0 97686 800 6 la_data_out[28]
port 291 nsew signal output
rlabel metal2 s 99194 0 99250 800 6 la_data_out[29]
port 292 nsew signal output
rlabel metal2 s 57794 0 57850 800 6 la_data_out[2]
port 293 nsew signal output
rlabel metal2 s 100666 0 100722 800 6 la_data_out[30]
port 294 nsew signal output
rlabel metal2 s 102230 0 102286 800 6 la_data_out[31]
port 295 nsew signal output
rlabel metal2 s 103794 0 103850 800 6 la_data_out[32]
port 296 nsew signal output
rlabel metal2 s 105266 0 105322 800 6 la_data_out[33]
port 297 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 la_data_out[34]
port 298 nsew signal output
rlabel metal2 s 108302 0 108358 800 6 la_data_out[35]
port 299 nsew signal output
rlabel metal2 s 109866 0 109922 800 6 la_data_out[36]
port 300 nsew signal output
rlabel metal2 s 111430 0 111486 800 6 la_data_out[37]
port 301 nsew signal output
rlabel metal2 s 112902 0 112958 800 6 la_data_out[38]
port 302 nsew signal output
rlabel metal2 s 114466 0 114522 800 6 la_data_out[39]
port 303 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 la_data_out[3]
port 304 nsew signal output
rlabel metal2 s 116030 0 116086 800 6 la_data_out[40]
port 305 nsew signal output
rlabel metal2 s 117502 0 117558 800 6 la_data_out[41]
port 306 nsew signal output
rlabel metal2 s 119066 0 119122 800 6 la_data_out[42]
port 307 nsew signal output
rlabel metal2 s 120630 0 120686 800 6 la_data_out[43]
port 308 nsew signal output
rlabel metal2 s 122102 0 122158 800 6 la_data_out[44]
port 309 nsew signal output
rlabel metal2 s 123666 0 123722 800 6 la_data_out[45]
port 310 nsew signal output
rlabel metal2 s 125230 0 125286 800 6 la_data_out[46]
port 311 nsew signal output
rlabel metal2 s 126702 0 126758 800 6 la_data_out[47]
port 312 nsew signal output
rlabel metal2 s 128266 0 128322 800 6 la_data_out[48]
port 313 nsew signal output
rlabel metal2 s 129738 0 129794 800 6 la_data_out[49]
port 314 nsew signal output
rlabel metal2 s 60922 0 60978 800 6 la_data_out[4]
port 315 nsew signal output
rlabel metal2 s 131302 0 131358 800 6 la_data_out[50]
port 316 nsew signal output
rlabel metal2 s 132866 0 132922 800 6 la_data_out[51]
port 317 nsew signal output
rlabel metal2 s 134338 0 134394 800 6 la_data_out[52]
port 318 nsew signal output
rlabel metal2 s 135902 0 135958 800 6 la_data_out[53]
port 319 nsew signal output
rlabel metal2 s 137466 0 137522 800 6 la_data_out[54]
port 320 nsew signal output
rlabel metal2 s 138938 0 138994 800 6 la_data_out[55]
port 321 nsew signal output
rlabel metal2 s 140502 0 140558 800 6 la_data_out[56]
port 322 nsew signal output
rlabel metal2 s 142066 0 142122 800 6 la_data_out[57]
port 323 nsew signal output
rlabel metal2 s 143538 0 143594 800 6 la_data_out[58]
port 324 nsew signal output
rlabel metal2 s 145102 0 145158 800 6 la_data_out[59]
port 325 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 la_data_out[5]
port 326 nsew signal output
rlabel metal2 s 146574 0 146630 800 6 la_data_out[60]
port 327 nsew signal output
rlabel metal2 s 148138 0 148194 800 6 la_data_out[61]
port 328 nsew signal output
rlabel metal2 s 149702 0 149758 800 6 la_data_out[62]
port 329 nsew signal output
rlabel metal2 s 151174 0 151230 800 6 la_data_out[63]
port 330 nsew signal output
rlabel metal2 s 152738 0 152794 800 6 la_data_out[64]
port 331 nsew signal output
rlabel metal2 s 154302 0 154358 800 6 la_data_out[65]
port 332 nsew signal output
rlabel metal2 s 155774 0 155830 800 6 la_data_out[66]
port 333 nsew signal output
rlabel metal2 s 157338 0 157394 800 6 la_data_out[67]
port 334 nsew signal output
rlabel metal2 s 158902 0 158958 800 6 la_data_out[68]
port 335 nsew signal output
rlabel metal2 s 160374 0 160430 800 6 la_data_out[69]
port 336 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 la_data_out[6]
port 337 nsew signal output
rlabel metal2 s 161938 0 161994 800 6 la_data_out[70]
port 338 nsew signal output
rlabel metal2 s 163502 0 163558 800 6 la_data_out[71]
port 339 nsew signal output
rlabel metal2 s 164974 0 165030 800 6 la_data_out[72]
port 340 nsew signal output
rlabel metal2 s 166538 0 166594 800 6 la_data_out[73]
port 341 nsew signal output
rlabel metal2 s 168010 0 168066 800 6 la_data_out[74]
port 342 nsew signal output
rlabel metal2 s 169574 0 169630 800 6 la_data_out[75]
port 343 nsew signal output
rlabel metal2 s 171138 0 171194 800 6 la_data_out[76]
port 344 nsew signal output
rlabel metal2 s 172610 0 172666 800 6 la_data_out[77]
port 345 nsew signal output
rlabel metal2 s 174174 0 174230 800 6 la_data_out[78]
port 346 nsew signal output
rlabel metal2 s 175738 0 175794 800 6 la_data_out[79]
port 347 nsew signal output
rlabel metal2 s 65522 0 65578 800 6 la_data_out[7]
port 348 nsew signal output
rlabel metal2 s 177210 0 177266 800 6 la_data_out[80]
port 349 nsew signal output
rlabel metal2 s 178774 0 178830 800 6 la_data_out[81]
port 350 nsew signal output
rlabel metal2 s 180338 0 180394 800 6 la_data_out[82]
port 351 nsew signal output
rlabel metal2 s 181810 0 181866 800 6 la_data_out[83]
port 352 nsew signal output
rlabel metal2 s 183374 0 183430 800 6 la_data_out[84]
port 353 nsew signal output
rlabel metal2 s 184846 0 184902 800 6 la_data_out[85]
port 354 nsew signal output
rlabel metal2 s 186410 0 186466 800 6 la_data_out[86]
port 355 nsew signal output
rlabel metal2 s 187974 0 188030 800 6 la_data_out[87]
port 356 nsew signal output
rlabel metal2 s 189446 0 189502 800 6 la_data_out[88]
port 357 nsew signal output
rlabel metal2 s 191010 0 191066 800 6 la_data_out[89]
port 358 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 la_data_out[8]
port 359 nsew signal output
rlabel metal2 s 192574 0 192630 800 6 la_data_out[90]
port 360 nsew signal output
rlabel metal2 s 194046 0 194102 800 6 la_data_out[91]
port 361 nsew signal output
rlabel metal2 s 195610 0 195666 800 6 la_data_out[92]
port 362 nsew signal output
rlabel metal2 s 197174 0 197230 800 6 la_data_out[93]
port 363 nsew signal output
rlabel metal2 s 198646 0 198702 800 6 la_data_out[94]
port 364 nsew signal output
rlabel metal2 s 200210 0 200266 800 6 la_data_out[95]
port 365 nsew signal output
rlabel metal2 s 201774 0 201830 800 6 la_data_out[96]
port 366 nsew signal output
rlabel metal2 s 203246 0 203302 800 6 la_data_out[97]
port 367 nsew signal output
rlabel metal2 s 204810 0 204866 800 6 la_data_out[98]
port 368 nsew signal output
rlabel metal2 s 206282 0 206338 800 6 la_data_out[99]
port 369 nsew signal output
rlabel metal2 s 68558 0 68614 800 6 la_data_out[9]
port 370 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 la_oen[0]
port 371 nsew signal input
rlabel metal2 s 208398 0 208454 800 6 la_oen[100]
port 372 nsew signal input
rlabel metal2 s 209870 0 209926 800 6 la_oen[101]
port 373 nsew signal input
rlabel metal2 s 211434 0 211490 800 6 la_oen[102]
port 374 nsew signal input
rlabel metal2 s 212998 0 213054 800 6 la_oen[103]
port 375 nsew signal input
rlabel metal2 s 214470 0 214526 800 6 la_oen[104]
port 376 nsew signal input
rlabel metal2 s 216034 0 216090 800 6 la_oen[105]
port 377 nsew signal input
rlabel metal2 s 217506 0 217562 800 6 la_oen[106]
port 378 nsew signal input
rlabel metal2 s 219070 0 219126 800 6 la_oen[107]
port 379 nsew signal input
rlabel metal2 s 220634 0 220690 800 6 la_oen[108]
port 380 nsew signal input
rlabel metal2 s 222106 0 222162 800 6 la_oen[109]
port 381 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 la_oen[10]
port 382 nsew signal input
rlabel metal2 s 223670 0 223726 800 6 la_oen[110]
port 383 nsew signal input
rlabel metal2 s 225234 0 225290 800 6 la_oen[111]
port 384 nsew signal input
rlabel metal2 s 226706 0 226762 800 6 la_oen[112]
port 385 nsew signal input
rlabel metal2 s 228270 0 228326 800 6 la_oen[113]
port 386 nsew signal input
rlabel metal2 s 229834 0 229890 800 6 la_oen[114]
port 387 nsew signal input
rlabel metal2 s 231306 0 231362 800 6 la_oen[115]
port 388 nsew signal input
rlabel metal2 s 232870 0 232926 800 6 la_oen[116]
port 389 nsew signal input
rlabel metal2 s 234434 0 234490 800 6 la_oen[117]
port 390 nsew signal input
rlabel metal2 s 235906 0 235962 800 6 la_oen[118]
port 391 nsew signal input
rlabel metal2 s 237470 0 237526 800 6 la_oen[119]
port 392 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 la_oen[11]
port 393 nsew signal input
rlabel metal2 s 238942 0 238998 800 6 la_oen[120]
port 394 nsew signal input
rlabel metal2 s 240506 0 240562 800 6 la_oen[121]
port 395 nsew signal input
rlabel metal2 s 242070 0 242126 800 6 la_oen[122]
port 396 nsew signal input
rlabel metal2 s 243542 0 243598 800 6 la_oen[123]
port 397 nsew signal input
rlabel metal2 s 245106 0 245162 800 6 la_oen[124]
port 398 nsew signal input
rlabel metal2 s 246670 0 246726 800 6 la_oen[125]
port 399 nsew signal input
rlabel metal2 s 248142 0 248198 800 6 la_oen[126]
port 400 nsew signal input
rlabel metal2 s 249706 0 249762 800 6 la_oen[127]
port 401 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_oen[12]
port 402 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 la_oen[13]
port 403 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 la_oen[14]
port 404 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_oen[15]
port 405 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_oen[16]
port 406 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_oen[17]
port 407 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_oen[18]
port 408 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_oen[19]
port 409 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_oen[1]
port 410 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_oen[20]
port 411 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_oen[21]
port 412 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_oen[22]
port 413 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 la_oen[23]
port 414 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_oen[24]
port 415 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_oen[25]
port 416 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 la_oen[26]
port 417 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_oen[27]
port 418 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 la_oen[28]
port 419 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 la_oen[29]
port 420 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 la_oen[2]
port 421 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 la_oen[30]
port 422 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 la_oen[31]
port 423 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 la_oen[32]
port 424 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_oen[33]
port 425 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 la_oen[34]
port 426 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 la_oen[35]
port 427 nsew signal input
rlabel metal2 s 110418 0 110474 800 6 la_oen[36]
port 428 nsew signal input
rlabel metal2 s 111890 0 111946 800 6 la_oen[37]
port 429 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 la_oen[38]
port 430 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 la_oen[39]
port 431 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_oen[3]
port 432 nsew signal input
rlabel metal2 s 116490 0 116546 800 6 la_oen[40]
port 433 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 la_oen[41]
port 434 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 la_oen[42]
port 435 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 la_oen[43]
port 436 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 la_oen[44]
port 437 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 la_oen[45]
port 438 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 la_oen[46]
port 439 nsew signal input
rlabel metal2 s 127254 0 127310 800 6 la_oen[47]
port 440 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 la_oen[48]
port 441 nsew signal input
rlabel metal2 s 130290 0 130346 800 6 la_oen[49]
port 442 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_oen[4]
port 443 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 la_oen[50]
port 444 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 la_oen[51]
port 445 nsew signal input
rlabel metal2 s 134890 0 134946 800 6 la_oen[52]
port 446 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 la_oen[53]
port 447 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 la_oen[54]
port 448 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 la_oen[55]
port 449 nsew signal input
rlabel metal2 s 140962 0 141018 800 6 la_oen[56]
port 450 nsew signal input
rlabel metal2 s 142526 0 142582 800 6 la_oen[57]
port 451 nsew signal input
rlabel metal2 s 144090 0 144146 800 6 la_oen[58]
port 452 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_oen[59]
port 453 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 la_oen[5]
port 454 nsew signal input
rlabel metal2 s 147126 0 147182 800 6 la_oen[60]
port 455 nsew signal input
rlabel metal2 s 148690 0 148746 800 6 la_oen[61]
port 456 nsew signal input
rlabel metal2 s 150162 0 150218 800 6 la_oen[62]
port 457 nsew signal input
rlabel metal2 s 151726 0 151782 800 6 la_oen[63]
port 458 nsew signal input
rlabel metal2 s 153290 0 153346 800 6 la_oen[64]
port 459 nsew signal input
rlabel metal2 s 154762 0 154818 800 6 la_oen[65]
port 460 nsew signal input
rlabel metal2 s 156326 0 156382 800 6 la_oen[66]
port 461 nsew signal input
rlabel metal2 s 157890 0 157946 800 6 la_oen[67]
port 462 nsew signal input
rlabel metal2 s 159362 0 159418 800 6 la_oen[68]
port 463 nsew signal input
rlabel metal2 s 160926 0 160982 800 6 la_oen[69]
port 464 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la_oen[6]
port 465 nsew signal input
rlabel metal2 s 162398 0 162454 800 6 la_oen[70]
port 466 nsew signal input
rlabel metal2 s 163962 0 164018 800 6 la_oen[71]
port 467 nsew signal input
rlabel metal2 s 165526 0 165582 800 6 la_oen[72]
port 468 nsew signal input
rlabel metal2 s 166998 0 167054 800 6 la_oen[73]
port 469 nsew signal input
rlabel metal2 s 168562 0 168618 800 6 la_oen[74]
port 470 nsew signal input
rlabel metal2 s 170126 0 170182 800 6 la_oen[75]
port 471 nsew signal input
rlabel metal2 s 171598 0 171654 800 6 la_oen[76]
port 472 nsew signal input
rlabel metal2 s 173162 0 173218 800 6 la_oen[77]
port 473 nsew signal input
rlabel metal2 s 174726 0 174782 800 6 la_oen[78]
port 474 nsew signal input
rlabel metal2 s 176198 0 176254 800 6 la_oen[79]
port 475 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_oen[7]
port 476 nsew signal input
rlabel metal2 s 177762 0 177818 800 6 la_oen[80]
port 477 nsew signal input
rlabel metal2 s 179234 0 179290 800 6 la_oen[81]
port 478 nsew signal input
rlabel metal2 s 180798 0 180854 800 6 la_oen[82]
port 479 nsew signal input
rlabel metal2 s 182362 0 182418 800 6 la_oen[83]
port 480 nsew signal input
rlabel metal2 s 183834 0 183890 800 6 la_oen[84]
port 481 nsew signal input
rlabel metal2 s 185398 0 185454 800 6 la_oen[85]
port 482 nsew signal input
rlabel metal2 s 186962 0 187018 800 6 la_oen[86]
port 483 nsew signal input
rlabel metal2 s 188434 0 188490 800 6 la_oen[87]
port 484 nsew signal input
rlabel metal2 s 189998 0 190054 800 6 la_oen[88]
port 485 nsew signal input
rlabel metal2 s 191562 0 191618 800 6 la_oen[89]
port 486 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_oen[8]
port 487 nsew signal input
rlabel metal2 s 193034 0 193090 800 6 la_oen[90]
port 488 nsew signal input
rlabel metal2 s 194598 0 194654 800 6 la_oen[91]
port 489 nsew signal input
rlabel metal2 s 196162 0 196218 800 6 la_oen[92]
port 490 nsew signal input
rlabel metal2 s 197634 0 197690 800 6 la_oen[93]
port 491 nsew signal input
rlabel metal2 s 199198 0 199254 800 6 la_oen[94]
port 492 nsew signal input
rlabel metal2 s 200670 0 200726 800 6 la_oen[95]
port 493 nsew signal input
rlabel metal2 s 202234 0 202290 800 6 la_oen[96]
port 494 nsew signal input
rlabel metal2 s 203798 0 203854 800 6 la_oen[97]
port 495 nsew signal input
rlabel metal2 s 205270 0 205326 800 6 la_oen[98]
port 496 nsew signal input
rlabel metal2 s 206834 0 206890 800 6 la_oen[99]
port 497 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 la_oen[9]
port 498 nsew signal input
rlabel metal4 s 4208 2128 4528 249744 6 vccd1
port 499 nsew power input
rlabel metal4 s 34928 2128 35248 249744 6 vccd1
port 499 nsew power input
rlabel metal4 s 65648 2128 65968 249744 6 vccd1
port 499 nsew power input
rlabel metal4 s 96368 2128 96688 249744 6 vccd1
port 499 nsew power input
rlabel metal4 s 127088 2128 127408 249744 6 vccd1
port 499 nsew power input
rlabel metal4 s 157808 2128 158128 249744 6 vccd1
port 499 nsew power input
rlabel metal4 s 188528 2128 188848 249744 6 vccd1
port 499 nsew power input
rlabel metal4 s 219248 2128 219568 249744 6 vccd1
port 499 nsew power input
rlabel metal4 s 19568 2128 19888 249744 6 vssd1
port 500 nsew ground input
rlabel metal4 s 50288 2128 50608 249744 6 vssd1
port 500 nsew ground input
rlabel metal4 s 81008 2128 81328 249744 6 vssd1
port 500 nsew ground input
rlabel metal4 s 111728 2128 112048 249744 6 vssd1
port 500 nsew ground input
rlabel metal4 s 142448 2128 142768 249744 6 vssd1
port 500 nsew ground input
rlabel metal4 s 173168 2128 173488 249744 6 vssd1
port 500 nsew ground input
rlabel metal4 s 203888 2128 204208 249744 6 vssd1
port 500 nsew ground input
rlabel metal4 s 234608 2128 234928 249744 6 vssd1
port 500 nsew ground input
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 501 nsew signal input
rlabel metal2 s 662 0 718 800 6 wb_rst_i
port 502 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 wbs_ack_o
port 503 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 wbs_adr_i[0]
port 504 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_adr_i[10]
port 505 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_adr_i[11]
port 506 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wbs_adr_i[12]
port 507 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_adr_i[13]
port 508 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_adr_i[14]
port 509 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 wbs_adr_i[15]
port 510 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_adr_i[16]
port 511 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 wbs_adr_i[17]
port 512 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 wbs_adr_i[18]
port 513 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 wbs_adr_i[19]
port 514 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_adr_i[1]
port 515 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_adr_i[20]
port 516 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 wbs_adr_i[21]
port 517 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 wbs_adr_i[22]
port 518 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wbs_adr_i[23]
port 519 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 wbs_adr_i[24]
port 520 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 wbs_adr_i[25]
port 521 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 wbs_adr_i[26]
port 522 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 wbs_adr_i[27]
port 523 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 wbs_adr_i[28]
port 524 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 wbs_adr_i[29]
port 525 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 wbs_adr_i[2]
port 526 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 wbs_adr_i[30]
port 527 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 wbs_adr_i[31]
port 528 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_adr_i[3]
port 529 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_adr_i[4]
port 530 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_adr_i[5]
port 531 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_adr_i[6]
port 532 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_adr_i[7]
port 533 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wbs_adr_i[8]
port 534 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_adr_i[9]
port 535 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_cyc_i
port 536 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_dat_i[0]
port 537 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_i[10]
port 538 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_dat_i[11]
port 539 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_dat_i[12]
port 540 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 wbs_dat_i[13]
port 541 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_i[14]
port 542 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_i[15]
port 543 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_i[16]
port 544 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 wbs_dat_i[17]
port 545 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wbs_dat_i[18]
port 546 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 wbs_dat_i[19]
port 547 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_dat_i[1]
port 548 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wbs_dat_i[20]
port 549 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 wbs_dat_i[21]
port 550 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 wbs_dat_i[22]
port 551 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 wbs_dat_i[23]
port 552 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_dat_i[24]
port 553 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 wbs_dat_i[25]
port 554 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 wbs_dat_i[26]
port 555 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 wbs_dat_i[27]
port 556 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 wbs_dat_i[28]
port 557 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 wbs_dat_i[29]
port 558 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_i[2]
port 559 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 wbs_dat_i[30]
port 560 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 wbs_dat_i[31]
port 561 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_i[3]
port 562 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_dat_i[4]
port 563 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_dat_i[5]
port 564 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_dat_i[6]
port 565 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_i[7]
port 566 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[8]
port 567 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_i[9]
port 568 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_dat_o[0]
port 569 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 wbs_dat_o[10]
port 570 nsew signal output
rlabel metal2 s 23110 0 23166 800 6 wbs_dat_o[11]
port 571 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_o[12]
port 572 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 wbs_dat_o[13]
port 573 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_o[14]
port 574 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 wbs_dat_o[15]
port 575 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 wbs_dat_o[16]
port 576 nsew signal output
rlabel metal2 s 32310 0 32366 800 6 wbs_dat_o[17]
port 577 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 wbs_dat_o[18]
port 578 nsew signal output
rlabel metal2 s 35346 0 35402 800 6 wbs_dat_o[19]
port 579 nsew signal output
rlabel metal2 s 6274 0 6330 800 6 wbs_dat_o[1]
port 580 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_o[20]
port 581 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 wbs_dat_o[21]
port 582 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 wbs_dat_o[22]
port 583 nsew signal output
rlabel metal2 s 41510 0 41566 800 6 wbs_dat_o[23]
port 584 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 wbs_dat_o[24]
port 585 nsew signal output
rlabel metal2 s 44546 0 44602 800 6 wbs_dat_o[25]
port 586 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 wbs_dat_o[26]
port 587 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 wbs_dat_o[27]
port 588 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 wbs_dat_o[28]
port 589 nsew signal output
rlabel metal2 s 50710 0 50766 800 6 wbs_dat_o[29]
port 590 nsew signal output
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_o[2]
port 591 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 wbs_dat_o[30]
port 592 nsew signal output
rlabel metal2 s 53746 0 53802 800 6 wbs_dat_o[31]
port 593 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_o[3]
port 594 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 wbs_dat_o[4]
port 595 nsew signal output
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_o[5]
port 596 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_o[6]
port 597 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 wbs_dat_o[7]
port 598 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 wbs_dat_o[8]
port 599 nsew signal output
rlabel metal2 s 20074 0 20130 800 6 wbs_dat_o[9]
port 600 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 wbs_sel_i[0]
port 601 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_sel_i[1]
port 602 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_sel_i[2]
port 603 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_sel_i[3]
port 604 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_stb_i
port 605 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_we_i
port 606 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 250060 252204
string LEFview TRUE
string GDS_FILE /project/openlane/accelerator_top/runs/accelerator_top/results/magic/accelerator_top.gds
string GDS_END 154770386
string GDS_START 1360094
<< end >>

