magic
tech sky130A
magscale 1 2
timestamp 1636397031
<< obsli1 >>
rect 1104 1377 278208 279089
<< obsm1 >>
rect 842 1368 278470 279120
<< metal2 >>
rect 1214 280659 1270 281459
rect 3606 280659 3662 281459
rect 6090 280659 6146 281459
rect 8482 280659 8538 281459
rect 10966 280659 11022 281459
rect 13450 280659 13506 281459
rect 15842 280659 15898 281459
rect 18326 280659 18382 281459
rect 20810 280659 20866 281459
rect 23202 280659 23258 281459
rect 25686 280659 25742 281459
rect 28078 280659 28134 281459
rect 30562 280659 30618 281459
rect 33046 280659 33102 281459
rect 35438 280659 35494 281459
rect 37922 280659 37978 281459
rect 40406 280659 40462 281459
rect 42798 280659 42854 281459
rect 45282 280659 45338 281459
rect 47766 280659 47822 281459
rect 50158 280659 50214 281459
rect 52642 280659 52698 281459
rect 55034 280659 55090 281459
rect 57518 280659 57574 281459
rect 60002 280659 60058 281459
rect 62394 280659 62450 281459
rect 64878 280659 64934 281459
rect 67362 280659 67418 281459
rect 69754 280659 69810 281459
rect 72238 280659 72294 281459
rect 74630 280659 74686 281459
rect 77114 280659 77170 281459
rect 79598 280659 79654 281459
rect 81990 280659 82046 281459
rect 84474 280659 84530 281459
rect 86958 280659 87014 281459
rect 89350 280659 89406 281459
rect 91834 280659 91890 281459
rect 94318 280659 94374 281459
rect 96710 280659 96766 281459
rect 99194 280659 99250 281459
rect 101586 280659 101642 281459
rect 104070 280659 104126 281459
rect 106554 280659 106610 281459
rect 108946 280659 109002 281459
rect 111430 280659 111486 281459
rect 113914 280659 113970 281459
rect 116306 280659 116362 281459
rect 118790 280659 118846 281459
rect 121182 280659 121238 281459
rect 123666 280659 123722 281459
rect 126150 280659 126206 281459
rect 128542 280659 128598 281459
rect 131026 280659 131082 281459
rect 133510 280659 133566 281459
rect 135902 280659 135958 281459
rect 138386 280659 138442 281459
rect 140870 280659 140926 281459
rect 143262 280659 143318 281459
rect 145746 280659 145802 281459
rect 148138 280659 148194 281459
rect 150622 280659 150678 281459
rect 153106 280659 153162 281459
rect 155498 280659 155554 281459
rect 157982 280659 158038 281459
rect 160466 280659 160522 281459
rect 162858 280659 162914 281459
rect 165342 280659 165398 281459
rect 167734 280659 167790 281459
rect 170218 280659 170274 281459
rect 172702 280659 172758 281459
rect 175094 280659 175150 281459
rect 177578 280659 177634 281459
rect 180062 280659 180118 281459
rect 182454 280659 182510 281459
rect 184938 280659 184994 281459
rect 187422 280659 187478 281459
rect 189814 280659 189870 281459
rect 192298 280659 192354 281459
rect 194690 280659 194746 281459
rect 197174 280659 197230 281459
rect 199658 280659 199714 281459
rect 202050 280659 202106 281459
rect 204534 280659 204590 281459
rect 207018 280659 207074 281459
rect 209410 280659 209466 281459
rect 211894 280659 211950 281459
rect 214286 280659 214342 281459
rect 216770 280659 216826 281459
rect 219254 280659 219310 281459
rect 221646 280659 221702 281459
rect 224130 280659 224186 281459
rect 226614 280659 226670 281459
rect 229006 280659 229062 281459
rect 231490 280659 231546 281459
rect 233974 280659 234030 281459
rect 236366 280659 236422 281459
rect 238850 280659 238906 281459
rect 241242 280659 241298 281459
rect 243726 280659 243782 281459
rect 246210 280659 246266 281459
rect 248602 280659 248658 281459
rect 251086 280659 251142 281459
rect 253570 280659 253626 281459
rect 255962 280659 256018 281459
rect 258446 280659 258502 281459
rect 260838 280659 260894 281459
rect 263322 280659 263378 281459
rect 265806 280659 265862 281459
rect 268198 280659 268254 281459
rect 270682 280659 270738 281459
rect 273166 280659 273222 281459
rect 275558 280659 275614 281459
rect 278042 280659 278098 281459
rect 294 0 350 800
rect 846 0 902 800
rect 1398 0 1454 800
rect 1950 0 2006 800
rect 2502 0 2558 800
rect 3054 0 3110 800
rect 3698 0 3754 800
rect 4250 0 4306 800
rect 4802 0 4858 800
rect 5354 0 5410 800
rect 5906 0 5962 800
rect 6550 0 6606 800
rect 7102 0 7158 800
rect 7654 0 7710 800
rect 8206 0 8262 800
rect 8758 0 8814 800
rect 9402 0 9458 800
rect 9954 0 10010 800
rect 10506 0 10562 800
rect 11058 0 11114 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12806 0 12862 800
rect 13358 0 13414 800
rect 13910 0 13966 800
rect 14462 0 14518 800
rect 15106 0 15162 800
rect 15658 0 15714 800
rect 16210 0 16266 800
rect 16762 0 16818 800
rect 17314 0 17370 800
rect 17958 0 18014 800
rect 18510 0 18566 800
rect 19062 0 19118 800
rect 19614 0 19670 800
rect 20166 0 20222 800
rect 20810 0 20866 800
rect 21362 0 21418 800
rect 21914 0 21970 800
rect 22466 0 22522 800
rect 23018 0 23074 800
rect 23662 0 23718 800
rect 24214 0 24270 800
rect 24766 0 24822 800
rect 25318 0 25374 800
rect 25870 0 25926 800
rect 26514 0 26570 800
rect 27066 0 27122 800
rect 27618 0 27674 800
rect 28170 0 28226 800
rect 28722 0 28778 800
rect 29274 0 29330 800
rect 29918 0 29974 800
rect 30470 0 30526 800
rect 31022 0 31078 800
rect 31574 0 31630 800
rect 32126 0 32182 800
rect 32770 0 32826 800
rect 33322 0 33378 800
rect 33874 0 33930 800
rect 34426 0 34482 800
rect 34978 0 35034 800
rect 35622 0 35678 800
rect 36174 0 36230 800
rect 36726 0 36782 800
rect 37278 0 37334 800
rect 37830 0 37886 800
rect 38474 0 38530 800
rect 39026 0 39082 800
rect 39578 0 39634 800
rect 40130 0 40186 800
rect 40682 0 40738 800
rect 41326 0 41382 800
rect 41878 0 41934 800
rect 42430 0 42486 800
rect 42982 0 43038 800
rect 43534 0 43590 800
rect 44178 0 44234 800
rect 44730 0 44786 800
rect 45282 0 45338 800
rect 45834 0 45890 800
rect 46386 0 46442 800
rect 47030 0 47086 800
rect 47582 0 47638 800
rect 48134 0 48190 800
rect 48686 0 48742 800
rect 49238 0 49294 800
rect 49882 0 49938 800
rect 50434 0 50490 800
rect 50986 0 51042 800
rect 51538 0 51594 800
rect 52090 0 52146 800
rect 52734 0 52790 800
rect 53286 0 53342 800
rect 53838 0 53894 800
rect 54390 0 54446 800
rect 54942 0 54998 800
rect 55586 0 55642 800
rect 56138 0 56194 800
rect 56690 0 56746 800
rect 57242 0 57298 800
rect 57794 0 57850 800
rect 58346 0 58402 800
rect 58990 0 59046 800
rect 59542 0 59598 800
rect 60094 0 60150 800
rect 60646 0 60702 800
rect 61198 0 61254 800
rect 61842 0 61898 800
rect 62394 0 62450 800
rect 62946 0 63002 800
rect 63498 0 63554 800
rect 64050 0 64106 800
rect 64694 0 64750 800
rect 65246 0 65302 800
rect 65798 0 65854 800
rect 66350 0 66406 800
rect 66902 0 66958 800
rect 67546 0 67602 800
rect 68098 0 68154 800
rect 68650 0 68706 800
rect 69202 0 69258 800
rect 69754 0 69810 800
rect 70398 0 70454 800
rect 70950 0 71006 800
rect 71502 0 71558 800
rect 72054 0 72110 800
rect 72606 0 72662 800
rect 73250 0 73306 800
rect 73802 0 73858 800
rect 74354 0 74410 800
rect 74906 0 74962 800
rect 75458 0 75514 800
rect 76102 0 76158 800
rect 76654 0 76710 800
rect 77206 0 77262 800
rect 77758 0 77814 800
rect 78310 0 78366 800
rect 78954 0 79010 800
rect 79506 0 79562 800
rect 80058 0 80114 800
rect 80610 0 80666 800
rect 81162 0 81218 800
rect 81806 0 81862 800
rect 82358 0 82414 800
rect 82910 0 82966 800
rect 83462 0 83518 800
rect 84014 0 84070 800
rect 84566 0 84622 800
rect 85210 0 85266 800
rect 85762 0 85818 800
rect 86314 0 86370 800
rect 86866 0 86922 800
rect 87418 0 87474 800
rect 88062 0 88118 800
rect 88614 0 88670 800
rect 89166 0 89222 800
rect 89718 0 89774 800
rect 90270 0 90326 800
rect 90914 0 90970 800
rect 91466 0 91522 800
rect 92018 0 92074 800
rect 92570 0 92626 800
rect 93122 0 93178 800
rect 93766 0 93822 800
rect 94318 0 94374 800
rect 94870 0 94926 800
rect 95422 0 95478 800
rect 95974 0 96030 800
rect 96618 0 96674 800
rect 97170 0 97226 800
rect 97722 0 97778 800
rect 98274 0 98330 800
rect 98826 0 98882 800
rect 99470 0 99526 800
rect 100022 0 100078 800
rect 100574 0 100630 800
rect 101126 0 101182 800
rect 101678 0 101734 800
rect 102322 0 102378 800
rect 102874 0 102930 800
rect 103426 0 103482 800
rect 103978 0 104034 800
rect 104530 0 104586 800
rect 105174 0 105230 800
rect 105726 0 105782 800
rect 106278 0 106334 800
rect 106830 0 106886 800
rect 107382 0 107438 800
rect 108026 0 108082 800
rect 108578 0 108634 800
rect 109130 0 109186 800
rect 109682 0 109738 800
rect 110234 0 110290 800
rect 110878 0 110934 800
rect 111430 0 111486 800
rect 111982 0 112038 800
rect 112534 0 112590 800
rect 113086 0 113142 800
rect 113638 0 113694 800
rect 114282 0 114338 800
rect 114834 0 114890 800
rect 115386 0 115442 800
rect 115938 0 115994 800
rect 116490 0 116546 800
rect 117134 0 117190 800
rect 117686 0 117742 800
rect 118238 0 118294 800
rect 118790 0 118846 800
rect 119342 0 119398 800
rect 119986 0 120042 800
rect 120538 0 120594 800
rect 121090 0 121146 800
rect 121642 0 121698 800
rect 122194 0 122250 800
rect 122838 0 122894 800
rect 123390 0 123446 800
rect 123942 0 123998 800
rect 124494 0 124550 800
rect 125046 0 125102 800
rect 125690 0 125746 800
rect 126242 0 126298 800
rect 126794 0 126850 800
rect 127346 0 127402 800
rect 127898 0 127954 800
rect 128542 0 128598 800
rect 129094 0 129150 800
rect 129646 0 129702 800
rect 130198 0 130254 800
rect 130750 0 130806 800
rect 131394 0 131450 800
rect 131946 0 132002 800
rect 132498 0 132554 800
rect 133050 0 133106 800
rect 133602 0 133658 800
rect 134246 0 134302 800
rect 134798 0 134854 800
rect 135350 0 135406 800
rect 135902 0 135958 800
rect 136454 0 136510 800
rect 137098 0 137154 800
rect 137650 0 137706 800
rect 138202 0 138258 800
rect 138754 0 138810 800
rect 139306 0 139362 800
rect 139950 0 140006 800
rect 140502 0 140558 800
rect 141054 0 141110 800
rect 141606 0 141662 800
rect 142158 0 142214 800
rect 142710 0 142766 800
rect 143354 0 143410 800
rect 143906 0 143962 800
rect 144458 0 144514 800
rect 145010 0 145066 800
rect 145562 0 145618 800
rect 146206 0 146262 800
rect 146758 0 146814 800
rect 147310 0 147366 800
rect 147862 0 147918 800
rect 148414 0 148470 800
rect 149058 0 149114 800
rect 149610 0 149666 800
rect 150162 0 150218 800
rect 150714 0 150770 800
rect 151266 0 151322 800
rect 151910 0 151966 800
rect 152462 0 152518 800
rect 153014 0 153070 800
rect 153566 0 153622 800
rect 154118 0 154174 800
rect 154762 0 154818 800
rect 155314 0 155370 800
rect 155866 0 155922 800
rect 156418 0 156474 800
rect 156970 0 157026 800
rect 157614 0 157670 800
rect 158166 0 158222 800
rect 158718 0 158774 800
rect 159270 0 159326 800
rect 159822 0 159878 800
rect 160466 0 160522 800
rect 161018 0 161074 800
rect 161570 0 161626 800
rect 162122 0 162178 800
rect 162674 0 162730 800
rect 163318 0 163374 800
rect 163870 0 163926 800
rect 164422 0 164478 800
rect 164974 0 165030 800
rect 165526 0 165582 800
rect 166170 0 166226 800
rect 166722 0 166778 800
rect 167274 0 167330 800
rect 167826 0 167882 800
rect 168378 0 168434 800
rect 168930 0 168986 800
rect 169574 0 169630 800
rect 170126 0 170182 800
rect 170678 0 170734 800
rect 171230 0 171286 800
rect 171782 0 171838 800
rect 172426 0 172482 800
rect 172978 0 173034 800
rect 173530 0 173586 800
rect 174082 0 174138 800
rect 174634 0 174690 800
rect 175278 0 175334 800
rect 175830 0 175886 800
rect 176382 0 176438 800
rect 176934 0 176990 800
rect 177486 0 177542 800
rect 178130 0 178186 800
rect 178682 0 178738 800
rect 179234 0 179290 800
rect 179786 0 179842 800
rect 180338 0 180394 800
rect 180982 0 181038 800
rect 181534 0 181590 800
rect 182086 0 182142 800
rect 182638 0 182694 800
rect 183190 0 183246 800
rect 183834 0 183890 800
rect 184386 0 184442 800
rect 184938 0 184994 800
rect 185490 0 185546 800
rect 186042 0 186098 800
rect 186686 0 186742 800
rect 187238 0 187294 800
rect 187790 0 187846 800
rect 188342 0 188398 800
rect 188894 0 188950 800
rect 189538 0 189594 800
rect 190090 0 190146 800
rect 190642 0 190698 800
rect 191194 0 191250 800
rect 191746 0 191802 800
rect 192390 0 192446 800
rect 192942 0 192998 800
rect 193494 0 193550 800
rect 194046 0 194102 800
rect 194598 0 194654 800
rect 195242 0 195298 800
rect 195794 0 195850 800
rect 196346 0 196402 800
rect 196898 0 196954 800
rect 197450 0 197506 800
rect 198002 0 198058 800
rect 198646 0 198702 800
rect 199198 0 199254 800
rect 199750 0 199806 800
rect 200302 0 200358 800
rect 200854 0 200910 800
rect 201498 0 201554 800
rect 202050 0 202106 800
rect 202602 0 202658 800
rect 203154 0 203210 800
rect 203706 0 203762 800
rect 204350 0 204406 800
rect 204902 0 204958 800
rect 205454 0 205510 800
rect 206006 0 206062 800
rect 206558 0 206614 800
rect 207202 0 207258 800
rect 207754 0 207810 800
rect 208306 0 208362 800
rect 208858 0 208914 800
rect 209410 0 209466 800
rect 210054 0 210110 800
rect 210606 0 210662 800
rect 211158 0 211214 800
rect 211710 0 211766 800
rect 212262 0 212318 800
rect 212906 0 212962 800
rect 213458 0 213514 800
rect 214010 0 214066 800
rect 214562 0 214618 800
rect 215114 0 215170 800
rect 215758 0 215814 800
rect 216310 0 216366 800
rect 216862 0 216918 800
rect 217414 0 217470 800
rect 217966 0 218022 800
rect 218610 0 218666 800
rect 219162 0 219218 800
rect 219714 0 219770 800
rect 220266 0 220322 800
rect 220818 0 220874 800
rect 221462 0 221518 800
rect 222014 0 222070 800
rect 222566 0 222622 800
rect 223118 0 223174 800
rect 223670 0 223726 800
rect 224222 0 224278 800
rect 224866 0 224922 800
rect 225418 0 225474 800
rect 225970 0 226026 800
rect 226522 0 226578 800
rect 227074 0 227130 800
rect 227718 0 227774 800
rect 228270 0 228326 800
rect 228822 0 228878 800
rect 229374 0 229430 800
rect 229926 0 229982 800
rect 230570 0 230626 800
rect 231122 0 231178 800
rect 231674 0 231730 800
rect 232226 0 232282 800
rect 232778 0 232834 800
rect 233422 0 233478 800
rect 233974 0 234030 800
rect 234526 0 234582 800
rect 235078 0 235134 800
rect 235630 0 235686 800
rect 236274 0 236330 800
rect 236826 0 236882 800
rect 237378 0 237434 800
rect 237930 0 237986 800
rect 238482 0 238538 800
rect 239126 0 239182 800
rect 239678 0 239734 800
rect 240230 0 240286 800
rect 240782 0 240838 800
rect 241334 0 241390 800
rect 241978 0 242034 800
rect 242530 0 242586 800
rect 243082 0 243138 800
rect 243634 0 243690 800
rect 244186 0 244242 800
rect 244830 0 244886 800
rect 245382 0 245438 800
rect 245934 0 245990 800
rect 246486 0 246542 800
rect 247038 0 247094 800
rect 247682 0 247738 800
rect 248234 0 248290 800
rect 248786 0 248842 800
rect 249338 0 249394 800
rect 249890 0 249946 800
rect 250534 0 250590 800
rect 251086 0 251142 800
rect 251638 0 251694 800
rect 252190 0 252246 800
rect 252742 0 252798 800
rect 253294 0 253350 800
rect 253938 0 253994 800
rect 254490 0 254546 800
rect 255042 0 255098 800
rect 255594 0 255650 800
rect 256146 0 256202 800
rect 256790 0 256846 800
rect 257342 0 257398 800
rect 257894 0 257950 800
rect 258446 0 258502 800
rect 258998 0 259054 800
rect 259642 0 259698 800
rect 260194 0 260250 800
rect 260746 0 260802 800
rect 261298 0 261354 800
rect 261850 0 261906 800
rect 262494 0 262550 800
rect 263046 0 263102 800
rect 263598 0 263654 800
rect 264150 0 264206 800
rect 264702 0 264758 800
rect 265346 0 265402 800
rect 265898 0 265954 800
rect 266450 0 266506 800
rect 267002 0 267058 800
rect 267554 0 267610 800
rect 268198 0 268254 800
rect 268750 0 268806 800
rect 269302 0 269358 800
rect 269854 0 269910 800
rect 270406 0 270462 800
rect 271050 0 271106 800
rect 271602 0 271658 800
rect 272154 0 272210 800
rect 272706 0 272762 800
rect 273258 0 273314 800
rect 273902 0 273958 800
rect 274454 0 274510 800
rect 275006 0 275062 800
rect 275558 0 275614 800
rect 276110 0 276166 800
rect 276754 0 276810 800
rect 277306 0 277362 800
rect 277858 0 277914 800
rect 278410 0 278466 800
rect 278962 0 279018 800
<< obsm2 >>
rect 294 280603 1158 280659
rect 1326 280603 3550 280659
rect 3718 280603 6034 280659
rect 6202 280603 8426 280659
rect 8594 280603 10910 280659
rect 11078 280603 13394 280659
rect 13562 280603 15786 280659
rect 15954 280603 18270 280659
rect 18438 280603 20754 280659
rect 20922 280603 23146 280659
rect 23314 280603 25630 280659
rect 25798 280603 28022 280659
rect 28190 280603 30506 280659
rect 30674 280603 32990 280659
rect 33158 280603 35382 280659
rect 35550 280603 37866 280659
rect 38034 280603 40350 280659
rect 40518 280603 42742 280659
rect 42910 280603 45226 280659
rect 45394 280603 47710 280659
rect 47878 280603 50102 280659
rect 50270 280603 52586 280659
rect 52754 280603 54978 280659
rect 55146 280603 57462 280659
rect 57630 280603 59946 280659
rect 60114 280603 62338 280659
rect 62506 280603 64822 280659
rect 64990 280603 67306 280659
rect 67474 280603 69698 280659
rect 69866 280603 72182 280659
rect 72350 280603 74574 280659
rect 74742 280603 77058 280659
rect 77226 280603 79542 280659
rect 79710 280603 81934 280659
rect 82102 280603 84418 280659
rect 84586 280603 86902 280659
rect 87070 280603 89294 280659
rect 89462 280603 91778 280659
rect 91946 280603 94262 280659
rect 94430 280603 96654 280659
rect 96822 280603 99138 280659
rect 99306 280603 101530 280659
rect 101698 280603 104014 280659
rect 104182 280603 106498 280659
rect 106666 280603 108890 280659
rect 109058 280603 111374 280659
rect 111542 280603 113858 280659
rect 114026 280603 116250 280659
rect 116418 280603 118734 280659
rect 118902 280603 121126 280659
rect 121294 280603 123610 280659
rect 123778 280603 126094 280659
rect 126262 280603 128486 280659
rect 128654 280603 130970 280659
rect 131138 280603 133454 280659
rect 133622 280603 135846 280659
rect 136014 280603 138330 280659
rect 138498 280603 140814 280659
rect 140982 280603 143206 280659
rect 143374 280603 145690 280659
rect 145858 280603 148082 280659
rect 148250 280603 150566 280659
rect 150734 280603 153050 280659
rect 153218 280603 155442 280659
rect 155610 280603 157926 280659
rect 158094 280603 160410 280659
rect 160578 280603 162802 280659
rect 162970 280603 165286 280659
rect 165454 280603 167678 280659
rect 167846 280603 170162 280659
rect 170330 280603 172646 280659
rect 172814 280603 175038 280659
rect 175206 280603 177522 280659
rect 177690 280603 180006 280659
rect 180174 280603 182398 280659
rect 182566 280603 184882 280659
rect 185050 280603 187366 280659
rect 187534 280603 189758 280659
rect 189926 280603 192242 280659
rect 192410 280603 194634 280659
rect 194802 280603 197118 280659
rect 197286 280603 199602 280659
rect 199770 280603 201994 280659
rect 202162 280603 204478 280659
rect 204646 280603 206962 280659
rect 207130 280603 209354 280659
rect 209522 280603 211838 280659
rect 212006 280603 214230 280659
rect 214398 280603 216714 280659
rect 216882 280603 219198 280659
rect 219366 280603 221590 280659
rect 221758 280603 224074 280659
rect 224242 280603 226558 280659
rect 226726 280603 228950 280659
rect 229118 280603 231434 280659
rect 231602 280603 233918 280659
rect 234086 280603 236310 280659
rect 236478 280603 238794 280659
rect 238962 280603 241186 280659
rect 241354 280603 243670 280659
rect 243838 280603 246154 280659
rect 246322 280603 248546 280659
rect 248714 280603 251030 280659
rect 251198 280603 253514 280659
rect 253682 280603 255906 280659
rect 256074 280603 258390 280659
rect 258558 280603 260782 280659
rect 260950 280603 263266 280659
rect 263434 280603 265750 280659
rect 265918 280603 268142 280659
rect 268310 280603 270626 280659
rect 270794 280603 273110 280659
rect 273278 280603 275502 280659
rect 275670 280603 277986 280659
rect 278154 280603 278464 280659
rect 294 856 278464 280603
rect 406 734 790 856
rect 958 734 1342 856
rect 1510 734 1894 856
rect 2062 734 2446 856
rect 2614 734 2998 856
rect 3166 734 3642 856
rect 3810 734 4194 856
rect 4362 734 4746 856
rect 4914 734 5298 856
rect 5466 734 5850 856
rect 6018 734 6494 856
rect 6662 734 7046 856
rect 7214 734 7598 856
rect 7766 734 8150 856
rect 8318 734 8702 856
rect 8870 734 9346 856
rect 9514 734 9898 856
rect 10066 734 10450 856
rect 10618 734 11002 856
rect 11170 734 11554 856
rect 11722 734 12198 856
rect 12366 734 12750 856
rect 12918 734 13302 856
rect 13470 734 13854 856
rect 14022 734 14406 856
rect 14574 734 15050 856
rect 15218 734 15602 856
rect 15770 734 16154 856
rect 16322 734 16706 856
rect 16874 734 17258 856
rect 17426 734 17902 856
rect 18070 734 18454 856
rect 18622 734 19006 856
rect 19174 734 19558 856
rect 19726 734 20110 856
rect 20278 734 20754 856
rect 20922 734 21306 856
rect 21474 734 21858 856
rect 22026 734 22410 856
rect 22578 734 22962 856
rect 23130 734 23606 856
rect 23774 734 24158 856
rect 24326 734 24710 856
rect 24878 734 25262 856
rect 25430 734 25814 856
rect 25982 734 26458 856
rect 26626 734 27010 856
rect 27178 734 27562 856
rect 27730 734 28114 856
rect 28282 734 28666 856
rect 28834 734 29218 856
rect 29386 734 29862 856
rect 30030 734 30414 856
rect 30582 734 30966 856
rect 31134 734 31518 856
rect 31686 734 32070 856
rect 32238 734 32714 856
rect 32882 734 33266 856
rect 33434 734 33818 856
rect 33986 734 34370 856
rect 34538 734 34922 856
rect 35090 734 35566 856
rect 35734 734 36118 856
rect 36286 734 36670 856
rect 36838 734 37222 856
rect 37390 734 37774 856
rect 37942 734 38418 856
rect 38586 734 38970 856
rect 39138 734 39522 856
rect 39690 734 40074 856
rect 40242 734 40626 856
rect 40794 734 41270 856
rect 41438 734 41822 856
rect 41990 734 42374 856
rect 42542 734 42926 856
rect 43094 734 43478 856
rect 43646 734 44122 856
rect 44290 734 44674 856
rect 44842 734 45226 856
rect 45394 734 45778 856
rect 45946 734 46330 856
rect 46498 734 46974 856
rect 47142 734 47526 856
rect 47694 734 48078 856
rect 48246 734 48630 856
rect 48798 734 49182 856
rect 49350 734 49826 856
rect 49994 734 50378 856
rect 50546 734 50930 856
rect 51098 734 51482 856
rect 51650 734 52034 856
rect 52202 734 52678 856
rect 52846 734 53230 856
rect 53398 734 53782 856
rect 53950 734 54334 856
rect 54502 734 54886 856
rect 55054 734 55530 856
rect 55698 734 56082 856
rect 56250 734 56634 856
rect 56802 734 57186 856
rect 57354 734 57738 856
rect 57906 734 58290 856
rect 58458 734 58934 856
rect 59102 734 59486 856
rect 59654 734 60038 856
rect 60206 734 60590 856
rect 60758 734 61142 856
rect 61310 734 61786 856
rect 61954 734 62338 856
rect 62506 734 62890 856
rect 63058 734 63442 856
rect 63610 734 63994 856
rect 64162 734 64638 856
rect 64806 734 65190 856
rect 65358 734 65742 856
rect 65910 734 66294 856
rect 66462 734 66846 856
rect 67014 734 67490 856
rect 67658 734 68042 856
rect 68210 734 68594 856
rect 68762 734 69146 856
rect 69314 734 69698 856
rect 69866 734 70342 856
rect 70510 734 70894 856
rect 71062 734 71446 856
rect 71614 734 71998 856
rect 72166 734 72550 856
rect 72718 734 73194 856
rect 73362 734 73746 856
rect 73914 734 74298 856
rect 74466 734 74850 856
rect 75018 734 75402 856
rect 75570 734 76046 856
rect 76214 734 76598 856
rect 76766 734 77150 856
rect 77318 734 77702 856
rect 77870 734 78254 856
rect 78422 734 78898 856
rect 79066 734 79450 856
rect 79618 734 80002 856
rect 80170 734 80554 856
rect 80722 734 81106 856
rect 81274 734 81750 856
rect 81918 734 82302 856
rect 82470 734 82854 856
rect 83022 734 83406 856
rect 83574 734 83958 856
rect 84126 734 84510 856
rect 84678 734 85154 856
rect 85322 734 85706 856
rect 85874 734 86258 856
rect 86426 734 86810 856
rect 86978 734 87362 856
rect 87530 734 88006 856
rect 88174 734 88558 856
rect 88726 734 89110 856
rect 89278 734 89662 856
rect 89830 734 90214 856
rect 90382 734 90858 856
rect 91026 734 91410 856
rect 91578 734 91962 856
rect 92130 734 92514 856
rect 92682 734 93066 856
rect 93234 734 93710 856
rect 93878 734 94262 856
rect 94430 734 94814 856
rect 94982 734 95366 856
rect 95534 734 95918 856
rect 96086 734 96562 856
rect 96730 734 97114 856
rect 97282 734 97666 856
rect 97834 734 98218 856
rect 98386 734 98770 856
rect 98938 734 99414 856
rect 99582 734 99966 856
rect 100134 734 100518 856
rect 100686 734 101070 856
rect 101238 734 101622 856
rect 101790 734 102266 856
rect 102434 734 102818 856
rect 102986 734 103370 856
rect 103538 734 103922 856
rect 104090 734 104474 856
rect 104642 734 105118 856
rect 105286 734 105670 856
rect 105838 734 106222 856
rect 106390 734 106774 856
rect 106942 734 107326 856
rect 107494 734 107970 856
rect 108138 734 108522 856
rect 108690 734 109074 856
rect 109242 734 109626 856
rect 109794 734 110178 856
rect 110346 734 110822 856
rect 110990 734 111374 856
rect 111542 734 111926 856
rect 112094 734 112478 856
rect 112646 734 113030 856
rect 113198 734 113582 856
rect 113750 734 114226 856
rect 114394 734 114778 856
rect 114946 734 115330 856
rect 115498 734 115882 856
rect 116050 734 116434 856
rect 116602 734 117078 856
rect 117246 734 117630 856
rect 117798 734 118182 856
rect 118350 734 118734 856
rect 118902 734 119286 856
rect 119454 734 119930 856
rect 120098 734 120482 856
rect 120650 734 121034 856
rect 121202 734 121586 856
rect 121754 734 122138 856
rect 122306 734 122782 856
rect 122950 734 123334 856
rect 123502 734 123886 856
rect 124054 734 124438 856
rect 124606 734 124990 856
rect 125158 734 125634 856
rect 125802 734 126186 856
rect 126354 734 126738 856
rect 126906 734 127290 856
rect 127458 734 127842 856
rect 128010 734 128486 856
rect 128654 734 129038 856
rect 129206 734 129590 856
rect 129758 734 130142 856
rect 130310 734 130694 856
rect 130862 734 131338 856
rect 131506 734 131890 856
rect 132058 734 132442 856
rect 132610 734 132994 856
rect 133162 734 133546 856
rect 133714 734 134190 856
rect 134358 734 134742 856
rect 134910 734 135294 856
rect 135462 734 135846 856
rect 136014 734 136398 856
rect 136566 734 137042 856
rect 137210 734 137594 856
rect 137762 734 138146 856
rect 138314 734 138698 856
rect 138866 734 139250 856
rect 139418 734 139894 856
rect 140062 734 140446 856
rect 140614 734 140998 856
rect 141166 734 141550 856
rect 141718 734 142102 856
rect 142270 734 142654 856
rect 142822 734 143298 856
rect 143466 734 143850 856
rect 144018 734 144402 856
rect 144570 734 144954 856
rect 145122 734 145506 856
rect 145674 734 146150 856
rect 146318 734 146702 856
rect 146870 734 147254 856
rect 147422 734 147806 856
rect 147974 734 148358 856
rect 148526 734 149002 856
rect 149170 734 149554 856
rect 149722 734 150106 856
rect 150274 734 150658 856
rect 150826 734 151210 856
rect 151378 734 151854 856
rect 152022 734 152406 856
rect 152574 734 152958 856
rect 153126 734 153510 856
rect 153678 734 154062 856
rect 154230 734 154706 856
rect 154874 734 155258 856
rect 155426 734 155810 856
rect 155978 734 156362 856
rect 156530 734 156914 856
rect 157082 734 157558 856
rect 157726 734 158110 856
rect 158278 734 158662 856
rect 158830 734 159214 856
rect 159382 734 159766 856
rect 159934 734 160410 856
rect 160578 734 160962 856
rect 161130 734 161514 856
rect 161682 734 162066 856
rect 162234 734 162618 856
rect 162786 734 163262 856
rect 163430 734 163814 856
rect 163982 734 164366 856
rect 164534 734 164918 856
rect 165086 734 165470 856
rect 165638 734 166114 856
rect 166282 734 166666 856
rect 166834 734 167218 856
rect 167386 734 167770 856
rect 167938 734 168322 856
rect 168490 734 168874 856
rect 169042 734 169518 856
rect 169686 734 170070 856
rect 170238 734 170622 856
rect 170790 734 171174 856
rect 171342 734 171726 856
rect 171894 734 172370 856
rect 172538 734 172922 856
rect 173090 734 173474 856
rect 173642 734 174026 856
rect 174194 734 174578 856
rect 174746 734 175222 856
rect 175390 734 175774 856
rect 175942 734 176326 856
rect 176494 734 176878 856
rect 177046 734 177430 856
rect 177598 734 178074 856
rect 178242 734 178626 856
rect 178794 734 179178 856
rect 179346 734 179730 856
rect 179898 734 180282 856
rect 180450 734 180926 856
rect 181094 734 181478 856
rect 181646 734 182030 856
rect 182198 734 182582 856
rect 182750 734 183134 856
rect 183302 734 183778 856
rect 183946 734 184330 856
rect 184498 734 184882 856
rect 185050 734 185434 856
rect 185602 734 185986 856
rect 186154 734 186630 856
rect 186798 734 187182 856
rect 187350 734 187734 856
rect 187902 734 188286 856
rect 188454 734 188838 856
rect 189006 734 189482 856
rect 189650 734 190034 856
rect 190202 734 190586 856
rect 190754 734 191138 856
rect 191306 734 191690 856
rect 191858 734 192334 856
rect 192502 734 192886 856
rect 193054 734 193438 856
rect 193606 734 193990 856
rect 194158 734 194542 856
rect 194710 734 195186 856
rect 195354 734 195738 856
rect 195906 734 196290 856
rect 196458 734 196842 856
rect 197010 734 197394 856
rect 197562 734 197946 856
rect 198114 734 198590 856
rect 198758 734 199142 856
rect 199310 734 199694 856
rect 199862 734 200246 856
rect 200414 734 200798 856
rect 200966 734 201442 856
rect 201610 734 201994 856
rect 202162 734 202546 856
rect 202714 734 203098 856
rect 203266 734 203650 856
rect 203818 734 204294 856
rect 204462 734 204846 856
rect 205014 734 205398 856
rect 205566 734 205950 856
rect 206118 734 206502 856
rect 206670 734 207146 856
rect 207314 734 207698 856
rect 207866 734 208250 856
rect 208418 734 208802 856
rect 208970 734 209354 856
rect 209522 734 209998 856
rect 210166 734 210550 856
rect 210718 734 211102 856
rect 211270 734 211654 856
rect 211822 734 212206 856
rect 212374 734 212850 856
rect 213018 734 213402 856
rect 213570 734 213954 856
rect 214122 734 214506 856
rect 214674 734 215058 856
rect 215226 734 215702 856
rect 215870 734 216254 856
rect 216422 734 216806 856
rect 216974 734 217358 856
rect 217526 734 217910 856
rect 218078 734 218554 856
rect 218722 734 219106 856
rect 219274 734 219658 856
rect 219826 734 220210 856
rect 220378 734 220762 856
rect 220930 734 221406 856
rect 221574 734 221958 856
rect 222126 734 222510 856
rect 222678 734 223062 856
rect 223230 734 223614 856
rect 223782 734 224166 856
rect 224334 734 224810 856
rect 224978 734 225362 856
rect 225530 734 225914 856
rect 226082 734 226466 856
rect 226634 734 227018 856
rect 227186 734 227662 856
rect 227830 734 228214 856
rect 228382 734 228766 856
rect 228934 734 229318 856
rect 229486 734 229870 856
rect 230038 734 230514 856
rect 230682 734 231066 856
rect 231234 734 231618 856
rect 231786 734 232170 856
rect 232338 734 232722 856
rect 232890 734 233366 856
rect 233534 734 233918 856
rect 234086 734 234470 856
rect 234638 734 235022 856
rect 235190 734 235574 856
rect 235742 734 236218 856
rect 236386 734 236770 856
rect 236938 734 237322 856
rect 237490 734 237874 856
rect 238042 734 238426 856
rect 238594 734 239070 856
rect 239238 734 239622 856
rect 239790 734 240174 856
rect 240342 734 240726 856
rect 240894 734 241278 856
rect 241446 734 241922 856
rect 242090 734 242474 856
rect 242642 734 243026 856
rect 243194 734 243578 856
rect 243746 734 244130 856
rect 244298 734 244774 856
rect 244942 734 245326 856
rect 245494 734 245878 856
rect 246046 734 246430 856
rect 246598 734 246982 856
rect 247150 734 247626 856
rect 247794 734 248178 856
rect 248346 734 248730 856
rect 248898 734 249282 856
rect 249450 734 249834 856
rect 250002 734 250478 856
rect 250646 734 251030 856
rect 251198 734 251582 856
rect 251750 734 252134 856
rect 252302 734 252686 856
rect 252854 734 253238 856
rect 253406 734 253882 856
rect 254050 734 254434 856
rect 254602 734 254986 856
rect 255154 734 255538 856
rect 255706 734 256090 856
rect 256258 734 256734 856
rect 256902 734 257286 856
rect 257454 734 257838 856
rect 258006 734 258390 856
rect 258558 734 258942 856
rect 259110 734 259586 856
rect 259754 734 260138 856
rect 260306 734 260690 856
rect 260858 734 261242 856
rect 261410 734 261794 856
rect 261962 734 262438 856
rect 262606 734 262990 856
rect 263158 734 263542 856
rect 263710 734 264094 856
rect 264262 734 264646 856
rect 264814 734 265290 856
rect 265458 734 265842 856
rect 266010 734 266394 856
rect 266562 734 266946 856
rect 267114 734 267498 856
rect 267666 734 268142 856
rect 268310 734 268694 856
rect 268862 734 269246 856
rect 269414 734 269798 856
rect 269966 734 270350 856
rect 270518 734 270994 856
rect 271162 734 271546 856
rect 271714 734 272098 856
rect 272266 734 272650 856
rect 272818 734 273202 856
rect 273370 734 273846 856
rect 274014 734 274398 856
rect 274566 734 274950 856
rect 275118 734 275502 856
rect 275670 734 276054 856
rect 276222 734 276698 856
rect 276866 734 277250 856
rect 277418 734 277802 856
rect 277970 734 278354 856
<< obsm3 >>
rect 289 1803 272307 279105
<< metal4 >>
rect 4208 2128 4528 279120
rect 19568 2128 19888 279120
rect 34928 2128 35248 279120
rect 50288 2128 50608 279120
rect 65648 2128 65968 279120
rect 81008 2128 81328 279120
rect 96368 2128 96688 279120
rect 111728 2128 112048 279120
rect 127088 2128 127408 279120
rect 142448 2128 142768 279120
rect 157808 2128 158128 279120
rect 173168 2128 173488 279120
rect 188528 2128 188848 279120
rect 203888 2128 204208 279120
rect 219248 2128 219568 279120
rect 234608 2128 234928 279120
rect 249968 2128 250288 279120
rect 265328 2128 265648 279120
<< obsm4 >>
rect 19195 25467 19488 240685
rect 19968 25467 34848 240685
rect 35328 25467 50208 240685
rect 50688 25467 65568 240685
rect 66048 25467 80928 240685
rect 81408 25467 96288 240685
rect 96768 25467 111648 240685
rect 112128 25467 127008 240685
rect 127488 25467 142368 240685
rect 142848 25467 157728 240685
rect 158208 25467 173088 240685
rect 173568 25467 188448 240685
rect 188928 25467 203808 240685
rect 204288 25467 219168 240685
rect 219648 25467 234528 240685
rect 235008 25467 249888 240685
rect 250368 25467 252941 240685
<< labels >>
rlabel metal2 s 1214 280659 1270 281459 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 74630 280659 74686 281459 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 81990 280659 82046 281459 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 89350 280659 89406 281459 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 96710 280659 96766 281459 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 104070 280659 104126 281459 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 111430 280659 111486 281459 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 118790 280659 118846 281459 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 126150 280659 126206 281459 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 133510 280659 133566 281459 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 140870 280659 140926 281459 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 8482 280659 8538 281459 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 148138 280659 148194 281459 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 155498 280659 155554 281459 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 162858 280659 162914 281459 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 170218 280659 170274 281459 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 177578 280659 177634 281459 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 184938 280659 184994 281459 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 192298 280659 192354 281459 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 199658 280659 199714 281459 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 207018 280659 207074 281459 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 214286 280659 214342 281459 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 15842 280659 15898 281459 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 221646 280659 221702 281459 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 229006 280659 229062 281459 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 236366 280659 236422 281459 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 243726 280659 243782 281459 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 251086 280659 251142 281459 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 258446 280659 258502 281459 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 265806 280659 265862 281459 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 273166 280659 273222 281459 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 23202 280659 23258 281459 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 30562 280659 30618 281459 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 37922 280659 37978 281459 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 45282 280659 45338 281459 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 52642 280659 52698 281459 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 60002 280659 60058 281459 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 67362 280659 67418 281459 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3606 280659 3662 281459 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 77114 280659 77170 281459 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 84474 280659 84530 281459 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 91834 280659 91890 281459 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 99194 280659 99250 281459 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 106554 280659 106610 281459 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 113914 280659 113970 281459 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 121182 280659 121238 281459 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 128542 280659 128598 281459 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 135902 280659 135958 281459 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 143262 280659 143318 281459 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 10966 280659 11022 281459 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 150622 280659 150678 281459 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 157982 280659 158038 281459 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 165342 280659 165398 281459 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 172702 280659 172758 281459 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 180062 280659 180118 281459 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 187422 280659 187478 281459 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 194690 280659 194746 281459 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 202050 280659 202106 281459 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 209410 280659 209466 281459 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 216770 280659 216826 281459 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 18326 280659 18382 281459 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 224130 280659 224186 281459 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 231490 280659 231546 281459 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 238850 280659 238906 281459 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 246210 280659 246266 281459 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 253570 280659 253626 281459 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 260838 280659 260894 281459 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 268198 280659 268254 281459 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 275558 280659 275614 281459 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 25686 280659 25742 281459 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 33046 280659 33102 281459 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 40406 280659 40462 281459 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 47766 280659 47822 281459 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 55034 280659 55090 281459 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 62394 280659 62450 281459 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 69754 280659 69810 281459 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 6090 280659 6146 281459 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 79598 280659 79654 281459 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 86958 280659 87014 281459 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 94318 280659 94374 281459 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 101586 280659 101642 281459 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 108946 280659 109002 281459 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 116306 280659 116362 281459 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 123666 280659 123722 281459 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 131026 280659 131082 281459 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 138386 280659 138442 281459 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 145746 280659 145802 281459 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 13450 280659 13506 281459 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 153106 280659 153162 281459 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 160466 280659 160522 281459 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 167734 280659 167790 281459 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 175094 280659 175150 281459 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 182454 280659 182510 281459 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 189814 280659 189870 281459 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 197174 280659 197230 281459 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 204534 280659 204590 281459 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 211894 280659 211950 281459 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 219254 280659 219310 281459 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 20810 280659 20866 281459 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 226614 280659 226670 281459 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 233974 280659 234030 281459 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 241242 280659 241298 281459 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 248602 280659 248658 281459 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 255962 280659 256018 281459 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 263322 280659 263378 281459 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 270682 280659 270738 281459 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 278042 280659 278098 281459 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 28078 280659 28134 281459 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 35438 280659 35494 281459 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 42798 280659 42854 281459 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 50158 280659 50214 281459 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 57518 280659 57574 281459 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 64878 280659 64934 281459 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 72238 280659 72294 281459 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 60646 0 60702 800 6 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 231674 0 231730 800 6 la_data_in[100]
port 116 nsew signal input
rlabel metal2 s 233422 0 233478 800 6 la_data_in[101]
port 117 nsew signal input
rlabel metal2 s 235078 0 235134 800 6 la_data_in[102]
port 118 nsew signal input
rlabel metal2 s 236826 0 236882 800 6 la_data_in[103]
port 119 nsew signal input
rlabel metal2 s 238482 0 238538 800 6 la_data_in[104]
port 120 nsew signal input
rlabel metal2 s 240230 0 240286 800 6 la_data_in[105]
port 121 nsew signal input
rlabel metal2 s 241978 0 242034 800 6 la_data_in[106]
port 122 nsew signal input
rlabel metal2 s 243634 0 243690 800 6 la_data_in[107]
port 123 nsew signal input
rlabel metal2 s 245382 0 245438 800 6 la_data_in[108]
port 124 nsew signal input
rlabel metal2 s 247038 0 247094 800 6 la_data_in[109]
port 125 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 la_data_in[10]
port 126 nsew signal input
rlabel metal2 s 248786 0 248842 800 6 la_data_in[110]
port 127 nsew signal input
rlabel metal2 s 250534 0 250590 800 6 la_data_in[111]
port 128 nsew signal input
rlabel metal2 s 252190 0 252246 800 6 la_data_in[112]
port 129 nsew signal input
rlabel metal2 s 253938 0 253994 800 6 la_data_in[113]
port 130 nsew signal input
rlabel metal2 s 255594 0 255650 800 6 la_data_in[114]
port 131 nsew signal input
rlabel metal2 s 257342 0 257398 800 6 la_data_in[115]
port 132 nsew signal input
rlabel metal2 s 258998 0 259054 800 6 la_data_in[116]
port 133 nsew signal input
rlabel metal2 s 260746 0 260802 800 6 la_data_in[117]
port 134 nsew signal input
rlabel metal2 s 262494 0 262550 800 6 la_data_in[118]
port 135 nsew signal input
rlabel metal2 s 264150 0 264206 800 6 la_data_in[119]
port 136 nsew signal input
rlabel metal2 s 79506 0 79562 800 6 la_data_in[11]
port 137 nsew signal input
rlabel metal2 s 265898 0 265954 800 6 la_data_in[120]
port 138 nsew signal input
rlabel metal2 s 267554 0 267610 800 6 la_data_in[121]
port 139 nsew signal input
rlabel metal2 s 269302 0 269358 800 6 la_data_in[122]
port 140 nsew signal input
rlabel metal2 s 271050 0 271106 800 6 la_data_in[123]
port 141 nsew signal input
rlabel metal2 s 272706 0 272762 800 6 la_data_in[124]
port 142 nsew signal input
rlabel metal2 s 274454 0 274510 800 6 la_data_in[125]
port 143 nsew signal input
rlabel metal2 s 276110 0 276166 800 6 la_data_in[126]
port 144 nsew signal input
rlabel metal2 s 277858 0 277914 800 6 la_data_in[127]
port 145 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_data_in[12]
port 146 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 la_data_in[13]
port 147 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 la_data_in[14]
port 148 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_data_in[15]
port 149 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_data_in[16]
port 150 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_data_in[17]
port 151 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 la_data_in[18]
port 152 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 la_data_in[19]
port 153 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 la_data_in[1]
port 154 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_data_in[20]
port 155 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_data_in[21]
port 156 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_data_in[22]
port 157 nsew signal input
rlabel metal2 s 100022 0 100078 800 6 la_data_in[23]
port 158 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_data_in[24]
port 159 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 la_data_in[25]
port 160 nsew signal input
rlabel metal2 s 105174 0 105230 800 6 la_data_in[26]
port 161 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 la_data_in[27]
port 162 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 la_data_in[28]
port 163 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 la_data_in[29]
port 164 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 la_data_in[2]
port 165 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 la_data_in[30]
port 166 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_data_in[31]
port 167 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 la_data_in[32]
port 168 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 la_data_in[33]
port 169 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 la_data_in[34]
port 170 nsew signal input
rlabel metal2 s 120538 0 120594 800 6 la_data_in[35]
port 171 nsew signal input
rlabel metal2 s 122194 0 122250 800 6 la_data_in[36]
port 172 nsew signal input
rlabel metal2 s 123942 0 123998 800 6 la_data_in[37]
port 173 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 la_data_in[38]
port 174 nsew signal input
rlabel metal2 s 127346 0 127402 800 6 la_data_in[39]
port 175 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 la_data_in[3]
port 176 nsew signal input
rlabel metal2 s 129094 0 129150 800 6 la_data_in[40]
port 177 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 la_data_in[41]
port 178 nsew signal input
rlabel metal2 s 132498 0 132554 800 6 la_data_in[42]
port 179 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 la_data_in[43]
port 180 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 la_data_in[44]
port 181 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 la_data_in[45]
port 182 nsew signal input
rlabel metal2 s 139306 0 139362 800 6 la_data_in[46]
port 183 nsew signal input
rlabel metal2 s 141054 0 141110 800 6 la_data_in[47]
port 184 nsew signal input
rlabel metal2 s 142710 0 142766 800 6 la_data_in[48]
port 185 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 la_data_in[49]
port 186 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_data_in[4]
port 187 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 la_data_in[50]
port 188 nsew signal input
rlabel metal2 s 147862 0 147918 800 6 la_data_in[51]
port 189 nsew signal input
rlabel metal2 s 149610 0 149666 800 6 la_data_in[52]
port 190 nsew signal input
rlabel metal2 s 151266 0 151322 800 6 la_data_in[53]
port 191 nsew signal input
rlabel metal2 s 153014 0 153070 800 6 la_data_in[54]
port 192 nsew signal input
rlabel metal2 s 154762 0 154818 800 6 la_data_in[55]
port 193 nsew signal input
rlabel metal2 s 156418 0 156474 800 6 la_data_in[56]
port 194 nsew signal input
rlabel metal2 s 158166 0 158222 800 6 la_data_in[57]
port 195 nsew signal input
rlabel metal2 s 159822 0 159878 800 6 la_data_in[58]
port 196 nsew signal input
rlabel metal2 s 161570 0 161626 800 6 la_data_in[59]
port 197 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_data_in[5]
port 198 nsew signal input
rlabel metal2 s 163318 0 163374 800 6 la_data_in[60]
port 199 nsew signal input
rlabel metal2 s 164974 0 165030 800 6 la_data_in[61]
port 200 nsew signal input
rlabel metal2 s 166722 0 166778 800 6 la_data_in[62]
port 201 nsew signal input
rlabel metal2 s 168378 0 168434 800 6 la_data_in[63]
port 202 nsew signal input
rlabel metal2 s 170126 0 170182 800 6 la_data_in[64]
port 203 nsew signal input
rlabel metal2 s 171782 0 171838 800 6 la_data_in[65]
port 204 nsew signal input
rlabel metal2 s 173530 0 173586 800 6 la_data_in[66]
port 205 nsew signal input
rlabel metal2 s 175278 0 175334 800 6 la_data_in[67]
port 206 nsew signal input
rlabel metal2 s 176934 0 176990 800 6 la_data_in[68]
port 207 nsew signal input
rlabel metal2 s 178682 0 178738 800 6 la_data_in[69]
port 208 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_data_in[6]
port 209 nsew signal input
rlabel metal2 s 180338 0 180394 800 6 la_data_in[70]
port 210 nsew signal input
rlabel metal2 s 182086 0 182142 800 6 la_data_in[71]
port 211 nsew signal input
rlabel metal2 s 183834 0 183890 800 6 la_data_in[72]
port 212 nsew signal input
rlabel metal2 s 185490 0 185546 800 6 la_data_in[73]
port 213 nsew signal input
rlabel metal2 s 187238 0 187294 800 6 la_data_in[74]
port 214 nsew signal input
rlabel metal2 s 188894 0 188950 800 6 la_data_in[75]
port 215 nsew signal input
rlabel metal2 s 190642 0 190698 800 6 la_data_in[76]
port 216 nsew signal input
rlabel metal2 s 192390 0 192446 800 6 la_data_in[77]
port 217 nsew signal input
rlabel metal2 s 194046 0 194102 800 6 la_data_in[78]
port 218 nsew signal input
rlabel metal2 s 195794 0 195850 800 6 la_data_in[79]
port 219 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 la_data_in[7]
port 220 nsew signal input
rlabel metal2 s 197450 0 197506 800 6 la_data_in[80]
port 221 nsew signal input
rlabel metal2 s 199198 0 199254 800 6 la_data_in[81]
port 222 nsew signal input
rlabel metal2 s 200854 0 200910 800 6 la_data_in[82]
port 223 nsew signal input
rlabel metal2 s 202602 0 202658 800 6 la_data_in[83]
port 224 nsew signal input
rlabel metal2 s 204350 0 204406 800 6 la_data_in[84]
port 225 nsew signal input
rlabel metal2 s 206006 0 206062 800 6 la_data_in[85]
port 226 nsew signal input
rlabel metal2 s 207754 0 207810 800 6 la_data_in[86]
port 227 nsew signal input
rlabel metal2 s 209410 0 209466 800 6 la_data_in[87]
port 228 nsew signal input
rlabel metal2 s 211158 0 211214 800 6 la_data_in[88]
port 229 nsew signal input
rlabel metal2 s 212906 0 212962 800 6 la_data_in[89]
port 230 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_data_in[8]
port 231 nsew signal input
rlabel metal2 s 214562 0 214618 800 6 la_data_in[90]
port 232 nsew signal input
rlabel metal2 s 216310 0 216366 800 6 la_data_in[91]
port 233 nsew signal input
rlabel metal2 s 217966 0 218022 800 6 la_data_in[92]
port 234 nsew signal input
rlabel metal2 s 219714 0 219770 800 6 la_data_in[93]
port 235 nsew signal input
rlabel metal2 s 221462 0 221518 800 6 la_data_in[94]
port 236 nsew signal input
rlabel metal2 s 223118 0 223174 800 6 la_data_in[95]
port 237 nsew signal input
rlabel metal2 s 224866 0 224922 800 6 la_data_in[96]
port 238 nsew signal input
rlabel metal2 s 226522 0 226578 800 6 la_data_in[97]
port 239 nsew signal input
rlabel metal2 s 228270 0 228326 800 6 la_data_in[98]
port 240 nsew signal input
rlabel metal2 s 229926 0 229982 800 6 la_data_in[99]
port 241 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 la_data_in[9]
port 242 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_data_out[0]
port 243 nsew signal output
rlabel metal2 s 232226 0 232282 800 6 la_data_out[100]
port 244 nsew signal output
rlabel metal2 s 233974 0 234030 800 6 la_data_out[101]
port 245 nsew signal output
rlabel metal2 s 235630 0 235686 800 6 la_data_out[102]
port 246 nsew signal output
rlabel metal2 s 237378 0 237434 800 6 la_data_out[103]
port 247 nsew signal output
rlabel metal2 s 239126 0 239182 800 6 la_data_out[104]
port 248 nsew signal output
rlabel metal2 s 240782 0 240838 800 6 la_data_out[105]
port 249 nsew signal output
rlabel metal2 s 242530 0 242586 800 6 la_data_out[106]
port 250 nsew signal output
rlabel metal2 s 244186 0 244242 800 6 la_data_out[107]
port 251 nsew signal output
rlabel metal2 s 245934 0 245990 800 6 la_data_out[108]
port 252 nsew signal output
rlabel metal2 s 247682 0 247738 800 6 la_data_out[109]
port 253 nsew signal output
rlabel metal2 s 78310 0 78366 800 6 la_data_out[10]
port 254 nsew signal output
rlabel metal2 s 249338 0 249394 800 6 la_data_out[110]
port 255 nsew signal output
rlabel metal2 s 251086 0 251142 800 6 la_data_out[111]
port 256 nsew signal output
rlabel metal2 s 252742 0 252798 800 6 la_data_out[112]
port 257 nsew signal output
rlabel metal2 s 254490 0 254546 800 6 la_data_out[113]
port 258 nsew signal output
rlabel metal2 s 256146 0 256202 800 6 la_data_out[114]
port 259 nsew signal output
rlabel metal2 s 257894 0 257950 800 6 la_data_out[115]
port 260 nsew signal output
rlabel metal2 s 259642 0 259698 800 6 la_data_out[116]
port 261 nsew signal output
rlabel metal2 s 261298 0 261354 800 6 la_data_out[117]
port 262 nsew signal output
rlabel metal2 s 263046 0 263102 800 6 la_data_out[118]
port 263 nsew signal output
rlabel metal2 s 264702 0 264758 800 6 la_data_out[119]
port 264 nsew signal output
rlabel metal2 s 80058 0 80114 800 6 la_data_out[11]
port 265 nsew signal output
rlabel metal2 s 266450 0 266506 800 6 la_data_out[120]
port 266 nsew signal output
rlabel metal2 s 268198 0 268254 800 6 la_data_out[121]
port 267 nsew signal output
rlabel metal2 s 269854 0 269910 800 6 la_data_out[122]
port 268 nsew signal output
rlabel metal2 s 271602 0 271658 800 6 la_data_out[123]
port 269 nsew signal output
rlabel metal2 s 273258 0 273314 800 6 la_data_out[124]
port 270 nsew signal output
rlabel metal2 s 275006 0 275062 800 6 la_data_out[125]
port 271 nsew signal output
rlabel metal2 s 276754 0 276810 800 6 la_data_out[126]
port 272 nsew signal output
rlabel metal2 s 278410 0 278466 800 6 la_data_out[127]
port 273 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 la_data_out[12]
port 274 nsew signal output
rlabel metal2 s 83462 0 83518 800 6 la_data_out[13]
port 275 nsew signal output
rlabel metal2 s 85210 0 85266 800 6 la_data_out[14]
port 276 nsew signal output
rlabel metal2 s 86866 0 86922 800 6 la_data_out[15]
port 277 nsew signal output
rlabel metal2 s 88614 0 88670 800 6 la_data_out[16]
port 278 nsew signal output
rlabel metal2 s 90270 0 90326 800 6 la_data_out[17]
port 279 nsew signal output
rlabel metal2 s 92018 0 92074 800 6 la_data_out[18]
port 280 nsew signal output
rlabel metal2 s 93766 0 93822 800 6 la_data_out[19]
port 281 nsew signal output
rlabel metal2 s 62946 0 63002 800 6 la_data_out[1]
port 282 nsew signal output
rlabel metal2 s 95422 0 95478 800 6 la_data_out[20]
port 283 nsew signal output
rlabel metal2 s 97170 0 97226 800 6 la_data_out[21]
port 284 nsew signal output
rlabel metal2 s 98826 0 98882 800 6 la_data_out[22]
port 285 nsew signal output
rlabel metal2 s 100574 0 100630 800 6 la_data_out[23]
port 286 nsew signal output
rlabel metal2 s 102322 0 102378 800 6 la_data_out[24]
port 287 nsew signal output
rlabel metal2 s 103978 0 104034 800 6 la_data_out[25]
port 288 nsew signal output
rlabel metal2 s 105726 0 105782 800 6 la_data_out[26]
port 289 nsew signal output
rlabel metal2 s 107382 0 107438 800 6 la_data_out[27]
port 290 nsew signal output
rlabel metal2 s 109130 0 109186 800 6 la_data_out[28]
port 291 nsew signal output
rlabel metal2 s 110878 0 110934 800 6 la_data_out[29]
port 292 nsew signal output
rlabel metal2 s 64694 0 64750 800 6 la_data_out[2]
port 293 nsew signal output
rlabel metal2 s 112534 0 112590 800 6 la_data_out[30]
port 294 nsew signal output
rlabel metal2 s 114282 0 114338 800 6 la_data_out[31]
port 295 nsew signal output
rlabel metal2 s 115938 0 115994 800 6 la_data_out[32]
port 296 nsew signal output
rlabel metal2 s 117686 0 117742 800 6 la_data_out[33]
port 297 nsew signal output
rlabel metal2 s 119342 0 119398 800 6 la_data_out[34]
port 298 nsew signal output
rlabel metal2 s 121090 0 121146 800 6 la_data_out[35]
port 299 nsew signal output
rlabel metal2 s 122838 0 122894 800 6 la_data_out[36]
port 300 nsew signal output
rlabel metal2 s 124494 0 124550 800 6 la_data_out[37]
port 301 nsew signal output
rlabel metal2 s 126242 0 126298 800 6 la_data_out[38]
port 302 nsew signal output
rlabel metal2 s 127898 0 127954 800 6 la_data_out[39]
port 303 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 la_data_out[3]
port 304 nsew signal output
rlabel metal2 s 129646 0 129702 800 6 la_data_out[40]
port 305 nsew signal output
rlabel metal2 s 131394 0 131450 800 6 la_data_out[41]
port 306 nsew signal output
rlabel metal2 s 133050 0 133106 800 6 la_data_out[42]
port 307 nsew signal output
rlabel metal2 s 134798 0 134854 800 6 la_data_out[43]
port 308 nsew signal output
rlabel metal2 s 136454 0 136510 800 6 la_data_out[44]
port 309 nsew signal output
rlabel metal2 s 138202 0 138258 800 6 la_data_out[45]
port 310 nsew signal output
rlabel metal2 s 139950 0 140006 800 6 la_data_out[46]
port 311 nsew signal output
rlabel metal2 s 141606 0 141662 800 6 la_data_out[47]
port 312 nsew signal output
rlabel metal2 s 143354 0 143410 800 6 la_data_out[48]
port 313 nsew signal output
rlabel metal2 s 145010 0 145066 800 6 la_data_out[49]
port 314 nsew signal output
rlabel metal2 s 68098 0 68154 800 6 la_data_out[4]
port 315 nsew signal output
rlabel metal2 s 146758 0 146814 800 6 la_data_out[50]
port 316 nsew signal output
rlabel metal2 s 148414 0 148470 800 6 la_data_out[51]
port 317 nsew signal output
rlabel metal2 s 150162 0 150218 800 6 la_data_out[52]
port 318 nsew signal output
rlabel metal2 s 151910 0 151966 800 6 la_data_out[53]
port 319 nsew signal output
rlabel metal2 s 153566 0 153622 800 6 la_data_out[54]
port 320 nsew signal output
rlabel metal2 s 155314 0 155370 800 6 la_data_out[55]
port 321 nsew signal output
rlabel metal2 s 156970 0 157026 800 6 la_data_out[56]
port 322 nsew signal output
rlabel metal2 s 158718 0 158774 800 6 la_data_out[57]
port 323 nsew signal output
rlabel metal2 s 160466 0 160522 800 6 la_data_out[58]
port 324 nsew signal output
rlabel metal2 s 162122 0 162178 800 6 la_data_out[59]
port 325 nsew signal output
rlabel metal2 s 69754 0 69810 800 6 la_data_out[5]
port 326 nsew signal output
rlabel metal2 s 163870 0 163926 800 6 la_data_out[60]
port 327 nsew signal output
rlabel metal2 s 165526 0 165582 800 6 la_data_out[61]
port 328 nsew signal output
rlabel metal2 s 167274 0 167330 800 6 la_data_out[62]
port 329 nsew signal output
rlabel metal2 s 168930 0 168986 800 6 la_data_out[63]
port 330 nsew signal output
rlabel metal2 s 170678 0 170734 800 6 la_data_out[64]
port 331 nsew signal output
rlabel metal2 s 172426 0 172482 800 6 la_data_out[65]
port 332 nsew signal output
rlabel metal2 s 174082 0 174138 800 6 la_data_out[66]
port 333 nsew signal output
rlabel metal2 s 175830 0 175886 800 6 la_data_out[67]
port 334 nsew signal output
rlabel metal2 s 177486 0 177542 800 6 la_data_out[68]
port 335 nsew signal output
rlabel metal2 s 179234 0 179290 800 6 la_data_out[69]
port 336 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 la_data_out[6]
port 337 nsew signal output
rlabel metal2 s 180982 0 181038 800 6 la_data_out[70]
port 338 nsew signal output
rlabel metal2 s 182638 0 182694 800 6 la_data_out[71]
port 339 nsew signal output
rlabel metal2 s 184386 0 184442 800 6 la_data_out[72]
port 340 nsew signal output
rlabel metal2 s 186042 0 186098 800 6 la_data_out[73]
port 341 nsew signal output
rlabel metal2 s 187790 0 187846 800 6 la_data_out[74]
port 342 nsew signal output
rlabel metal2 s 189538 0 189594 800 6 la_data_out[75]
port 343 nsew signal output
rlabel metal2 s 191194 0 191250 800 6 la_data_out[76]
port 344 nsew signal output
rlabel metal2 s 192942 0 192998 800 6 la_data_out[77]
port 345 nsew signal output
rlabel metal2 s 194598 0 194654 800 6 la_data_out[78]
port 346 nsew signal output
rlabel metal2 s 196346 0 196402 800 6 la_data_out[79]
port 347 nsew signal output
rlabel metal2 s 73250 0 73306 800 6 la_data_out[7]
port 348 nsew signal output
rlabel metal2 s 198002 0 198058 800 6 la_data_out[80]
port 349 nsew signal output
rlabel metal2 s 199750 0 199806 800 6 la_data_out[81]
port 350 nsew signal output
rlabel metal2 s 201498 0 201554 800 6 la_data_out[82]
port 351 nsew signal output
rlabel metal2 s 203154 0 203210 800 6 la_data_out[83]
port 352 nsew signal output
rlabel metal2 s 204902 0 204958 800 6 la_data_out[84]
port 353 nsew signal output
rlabel metal2 s 206558 0 206614 800 6 la_data_out[85]
port 354 nsew signal output
rlabel metal2 s 208306 0 208362 800 6 la_data_out[86]
port 355 nsew signal output
rlabel metal2 s 210054 0 210110 800 6 la_data_out[87]
port 356 nsew signal output
rlabel metal2 s 211710 0 211766 800 6 la_data_out[88]
port 357 nsew signal output
rlabel metal2 s 213458 0 213514 800 6 la_data_out[89]
port 358 nsew signal output
rlabel metal2 s 74906 0 74962 800 6 la_data_out[8]
port 359 nsew signal output
rlabel metal2 s 215114 0 215170 800 6 la_data_out[90]
port 360 nsew signal output
rlabel metal2 s 216862 0 216918 800 6 la_data_out[91]
port 361 nsew signal output
rlabel metal2 s 218610 0 218666 800 6 la_data_out[92]
port 362 nsew signal output
rlabel metal2 s 220266 0 220322 800 6 la_data_out[93]
port 363 nsew signal output
rlabel metal2 s 222014 0 222070 800 6 la_data_out[94]
port 364 nsew signal output
rlabel metal2 s 223670 0 223726 800 6 la_data_out[95]
port 365 nsew signal output
rlabel metal2 s 225418 0 225474 800 6 la_data_out[96]
port 366 nsew signal output
rlabel metal2 s 227074 0 227130 800 6 la_data_out[97]
port 367 nsew signal output
rlabel metal2 s 228822 0 228878 800 6 la_data_out[98]
port 368 nsew signal output
rlabel metal2 s 230570 0 230626 800 6 la_data_out[99]
port 369 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 la_data_out[9]
port 370 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 la_oen[0]
port 371 nsew signal input
rlabel metal2 s 232778 0 232834 800 6 la_oen[100]
port 372 nsew signal input
rlabel metal2 s 234526 0 234582 800 6 la_oen[101]
port 373 nsew signal input
rlabel metal2 s 236274 0 236330 800 6 la_oen[102]
port 374 nsew signal input
rlabel metal2 s 237930 0 237986 800 6 la_oen[103]
port 375 nsew signal input
rlabel metal2 s 239678 0 239734 800 6 la_oen[104]
port 376 nsew signal input
rlabel metal2 s 241334 0 241390 800 6 la_oen[105]
port 377 nsew signal input
rlabel metal2 s 243082 0 243138 800 6 la_oen[106]
port 378 nsew signal input
rlabel metal2 s 244830 0 244886 800 6 la_oen[107]
port 379 nsew signal input
rlabel metal2 s 246486 0 246542 800 6 la_oen[108]
port 380 nsew signal input
rlabel metal2 s 248234 0 248290 800 6 la_oen[109]
port 381 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_oen[10]
port 382 nsew signal input
rlabel metal2 s 249890 0 249946 800 6 la_oen[110]
port 383 nsew signal input
rlabel metal2 s 251638 0 251694 800 6 la_oen[111]
port 384 nsew signal input
rlabel metal2 s 253294 0 253350 800 6 la_oen[112]
port 385 nsew signal input
rlabel metal2 s 255042 0 255098 800 6 la_oen[113]
port 386 nsew signal input
rlabel metal2 s 256790 0 256846 800 6 la_oen[114]
port 387 nsew signal input
rlabel metal2 s 258446 0 258502 800 6 la_oen[115]
port 388 nsew signal input
rlabel metal2 s 260194 0 260250 800 6 la_oen[116]
port 389 nsew signal input
rlabel metal2 s 261850 0 261906 800 6 la_oen[117]
port 390 nsew signal input
rlabel metal2 s 263598 0 263654 800 6 la_oen[118]
port 391 nsew signal input
rlabel metal2 s 265346 0 265402 800 6 la_oen[119]
port 392 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 la_oen[11]
port 393 nsew signal input
rlabel metal2 s 267002 0 267058 800 6 la_oen[120]
port 394 nsew signal input
rlabel metal2 s 268750 0 268806 800 6 la_oen[121]
port 395 nsew signal input
rlabel metal2 s 270406 0 270462 800 6 la_oen[122]
port 396 nsew signal input
rlabel metal2 s 272154 0 272210 800 6 la_oen[123]
port 397 nsew signal input
rlabel metal2 s 273902 0 273958 800 6 la_oen[124]
port 398 nsew signal input
rlabel metal2 s 275558 0 275614 800 6 la_oen[125]
port 399 nsew signal input
rlabel metal2 s 277306 0 277362 800 6 la_oen[126]
port 400 nsew signal input
rlabel metal2 s 278962 0 279018 800 6 la_oen[127]
port 401 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_oen[12]
port 402 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_oen[13]
port 403 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_oen[14]
port 404 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_oen[15]
port 405 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_oen[16]
port 406 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_oen[17]
port 407 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_oen[18]
port 408 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 la_oen[19]
port 409 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_oen[1]
port 410 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_oen[20]
port 411 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 la_oen[21]
port 412 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_oen[22]
port 413 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_oen[23]
port 414 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 la_oen[24]
port 415 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 la_oen[25]
port 416 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 la_oen[26]
port 417 nsew signal input
rlabel metal2 s 108026 0 108082 800 6 la_oen[27]
port 418 nsew signal input
rlabel metal2 s 109682 0 109738 800 6 la_oen[28]
port 419 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 la_oen[29]
port 420 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 la_oen[2]
port 421 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 la_oen[30]
port 422 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 la_oen[31]
port 423 nsew signal input
rlabel metal2 s 116490 0 116546 800 6 la_oen[32]
port 424 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 la_oen[33]
port 425 nsew signal input
rlabel metal2 s 119986 0 120042 800 6 la_oen[34]
port 426 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 la_oen[35]
port 427 nsew signal input
rlabel metal2 s 123390 0 123446 800 6 la_oen[36]
port 428 nsew signal input
rlabel metal2 s 125046 0 125102 800 6 la_oen[37]
port 429 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 la_oen[38]
port 430 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 la_oen[39]
port 431 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 la_oen[3]
port 432 nsew signal input
rlabel metal2 s 130198 0 130254 800 6 la_oen[40]
port 433 nsew signal input
rlabel metal2 s 131946 0 132002 800 6 la_oen[41]
port 434 nsew signal input
rlabel metal2 s 133602 0 133658 800 6 la_oen[42]
port 435 nsew signal input
rlabel metal2 s 135350 0 135406 800 6 la_oen[43]
port 436 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 la_oen[44]
port 437 nsew signal input
rlabel metal2 s 138754 0 138810 800 6 la_oen[45]
port 438 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 la_oen[46]
port 439 nsew signal input
rlabel metal2 s 142158 0 142214 800 6 la_oen[47]
port 440 nsew signal input
rlabel metal2 s 143906 0 143962 800 6 la_oen[48]
port 441 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_oen[49]
port 442 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 la_oen[4]
port 443 nsew signal input
rlabel metal2 s 147310 0 147366 800 6 la_oen[50]
port 444 nsew signal input
rlabel metal2 s 149058 0 149114 800 6 la_oen[51]
port 445 nsew signal input
rlabel metal2 s 150714 0 150770 800 6 la_oen[52]
port 446 nsew signal input
rlabel metal2 s 152462 0 152518 800 6 la_oen[53]
port 447 nsew signal input
rlabel metal2 s 154118 0 154174 800 6 la_oen[54]
port 448 nsew signal input
rlabel metal2 s 155866 0 155922 800 6 la_oen[55]
port 449 nsew signal input
rlabel metal2 s 157614 0 157670 800 6 la_oen[56]
port 450 nsew signal input
rlabel metal2 s 159270 0 159326 800 6 la_oen[57]
port 451 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 la_oen[58]
port 452 nsew signal input
rlabel metal2 s 162674 0 162730 800 6 la_oen[59]
port 453 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_oen[5]
port 454 nsew signal input
rlabel metal2 s 164422 0 164478 800 6 la_oen[60]
port 455 nsew signal input
rlabel metal2 s 166170 0 166226 800 6 la_oen[61]
port 456 nsew signal input
rlabel metal2 s 167826 0 167882 800 6 la_oen[62]
port 457 nsew signal input
rlabel metal2 s 169574 0 169630 800 6 la_oen[63]
port 458 nsew signal input
rlabel metal2 s 171230 0 171286 800 6 la_oen[64]
port 459 nsew signal input
rlabel metal2 s 172978 0 173034 800 6 la_oen[65]
port 460 nsew signal input
rlabel metal2 s 174634 0 174690 800 6 la_oen[66]
port 461 nsew signal input
rlabel metal2 s 176382 0 176438 800 6 la_oen[67]
port 462 nsew signal input
rlabel metal2 s 178130 0 178186 800 6 la_oen[68]
port 463 nsew signal input
rlabel metal2 s 179786 0 179842 800 6 la_oen[69]
port 464 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_oen[6]
port 465 nsew signal input
rlabel metal2 s 181534 0 181590 800 6 la_oen[70]
port 466 nsew signal input
rlabel metal2 s 183190 0 183246 800 6 la_oen[71]
port 467 nsew signal input
rlabel metal2 s 184938 0 184994 800 6 la_oen[72]
port 468 nsew signal input
rlabel metal2 s 186686 0 186742 800 6 la_oen[73]
port 469 nsew signal input
rlabel metal2 s 188342 0 188398 800 6 la_oen[74]
port 470 nsew signal input
rlabel metal2 s 190090 0 190146 800 6 la_oen[75]
port 471 nsew signal input
rlabel metal2 s 191746 0 191802 800 6 la_oen[76]
port 472 nsew signal input
rlabel metal2 s 193494 0 193550 800 6 la_oen[77]
port 473 nsew signal input
rlabel metal2 s 195242 0 195298 800 6 la_oen[78]
port 474 nsew signal input
rlabel metal2 s 196898 0 196954 800 6 la_oen[79]
port 475 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_oen[7]
port 476 nsew signal input
rlabel metal2 s 198646 0 198702 800 6 la_oen[80]
port 477 nsew signal input
rlabel metal2 s 200302 0 200358 800 6 la_oen[81]
port 478 nsew signal input
rlabel metal2 s 202050 0 202106 800 6 la_oen[82]
port 479 nsew signal input
rlabel metal2 s 203706 0 203762 800 6 la_oen[83]
port 480 nsew signal input
rlabel metal2 s 205454 0 205510 800 6 la_oen[84]
port 481 nsew signal input
rlabel metal2 s 207202 0 207258 800 6 la_oen[85]
port 482 nsew signal input
rlabel metal2 s 208858 0 208914 800 6 la_oen[86]
port 483 nsew signal input
rlabel metal2 s 210606 0 210662 800 6 la_oen[87]
port 484 nsew signal input
rlabel metal2 s 212262 0 212318 800 6 la_oen[88]
port 485 nsew signal input
rlabel metal2 s 214010 0 214066 800 6 la_oen[89]
port 486 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_oen[8]
port 487 nsew signal input
rlabel metal2 s 215758 0 215814 800 6 la_oen[90]
port 488 nsew signal input
rlabel metal2 s 217414 0 217470 800 6 la_oen[91]
port 489 nsew signal input
rlabel metal2 s 219162 0 219218 800 6 la_oen[92]
port 490 nsew signal input
rlabel metal2 s 220818 0 220874 800 6 la_oen[93]
port 491 nsew signal input
rlabel metal2 s 222566 0 222622 800 6 la_oen[94]
port 492 nsew signal input
rlabel metal2 s 224222 0 224278 800 6 la_oen[95]
port 493 nsew signal input
rlabel metal2 s 225970 0 226026 800 6 la_oen[96]
port 494 nsew signal input
rlabel metal2 s 227718 0 227774 800 6 la_oen[97]
port 495 nsew signal input
rlabel metal2 s 229374 0 229430 800 6 la_oen[98]
port 496 nsew signal input
rlabel metal2 s 231122 0 231178 800 6 la_oen[99]
port 497 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_oen[9]
port 498 nsew signal input
rlabel metal4 s 4208 2128 4528 279120 6 vccd1
port 499 nsew power input
rlabel metal4 s 34928 2128 35248 279120 6 vccd1
port 499 nsew power input
rlabel metal4 s 65648 2128 65968 279120 6 vccd1
port 499 nsew power input
rlabel metal4 s 96368 2128 96688 279120 6 vccd1
port 499 nsew power input
rlabel metal4 s 127088 2128 127408 279120 6 vccd1
port 499 nsew power input
rlabel metal4 s 157808 2128 158128 279120 6 vccd1
port 499 nsew power input
rlabel metal4 s 188528 2128 188848 279120 6 vccd1
port 499 nsew power input
rlabel metal4 s 219248 2128 219568 279120 6 vccd1
port 499 nsew power input
rlabel metal4 s 249968 2128 250288 279120 6 vccd1
port 499 nsew power input
rlabel metal4 s 19568 2128 19888 279120 6 vssd1
port 500 nsew ground input
rlabel metal4 s 50288 2128 50608 279120 6 vssd1
port 500 nsew ground input
rlabel metal4 s 81008 2128 81328 279120 6 vssd1
port 500 nsew ground input
rlabel metal4 s 111728 2128 112048 279120 6 vssd1
port 500 nsew ground input
rlabel metal4 s 142448 2128 142768 279120 6 vssd1
port 500 nsew ground input
rlabel metal4 s 173168 2128 173488 279120 6 vssd1
port 500 nsew ground input
rlabel metal4 s 203888 2128 204208 279120 6 vssd1
port 500 nsew ground input
rlabel metal4 s 234608 2128 234928 279120 6 vssd1
port 500 nsew ground input
rlabel metal4 s 265328 2128 265648 279120 6 vssd1
port 500 nsew ground input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 501 nsew signal input
rlabel metal2 s 846 0 902 800 6 wb_rst_i
port 502 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_ack_o
port 503 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[0]
port 504 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_adr_i[10]
port 505 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_adr_i[11]
port 506 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 wbs_adr_i[12]
port 507 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 wbs_adr_i[13]
port 508 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_adr_i[14]
port 509 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_adr_i[15]
port 510 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wbs_adr_i[16]
port 511 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 wbs_adr_i[17]
port 512 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 wbs_adr_i[18]
port 513 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 wbs_adr_i[19]
port 514 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_adr_i[1]
port 515 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 wbs_adr_i[20]
port 516 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 wbs_adr_i[21]
port 517 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 wbs_adr_i[22]
port 518 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 wbs_adr_i[23]
port 519 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 wbs_adr_i[24]
port 520 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 wbs_adr_i[25]
port 521 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 wbs_adr_i[26]
port 522 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 wbs_adr_i[27]
port 523 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 wbs_adr_i[28]
port 524 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 wbs_adr_i[29]
port 525 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[2]
port 526 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 wbs_adr_i[30]
port 527 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 wbs_adr_i[31]
port 528 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 wbs_adr_i[3]
port 529 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_adr_i[4]
port 530 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_adr_i[5]
port 531 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 wbs_adr_i[6]
port 532 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[7]
port 533 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 wbs_adr_i[8]
port 534 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_adr_i[9]
port 535 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_cyc_i
port 536 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_dat_i[0]
port 537 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wbs_dat_i[10]
port 538 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_dat_i[11]
port 539 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 wbs_dat_i[12]
port 540 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_i[13]
port 541 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_i[14]
port 542 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_i[15]
port 543 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wbs_dat_i[16]
port 544 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 wbs_dat_i[17]
port 545 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 wbs_dat_i[18]
port 546 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 wbs_dat_i[19]
port 547 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_i[1]
port 548 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 wbs_dat_i[20]
port 549 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 wbs_dat_i[21]
port 550 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 wbs_dat_i[22]
port 551 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 wbs_dat_i[23]
port 552 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 wbs_dat_i[24]
port 553 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 wbs_dat_i[25]
port 554 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 wbs_dat_i[26]
port 555 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 wbs_dat_i[27]
port 556 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 wbs_dat_i[28]
port 557 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 wbs_dat_i[29]
port 558 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_i[2]
port 559 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 wbs_dat_i[30]
port 560 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 wbs_dat_i[31]
port 561 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_i[3]
port 562 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_dat_i[4]
port 563 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_i[5]
port 564 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_dat_i[6]
port 565 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wbs_dat_i[7]
port 566 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_i[8]
port 567 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wbs_dat_i[9]
port 568 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_dat_o[0]
port 569 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 wbs_dat_o[10]
port 570 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 wbs_dat_o[11]
port 571 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 wbs_dat_o[12]
port 572 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 wbs_dat_o[13]
port 573 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 wbs_dat_o[14]
port 574 nsew signal output
rlabel metal2 s 32770 0 32826 800 6 wbs_dat_o[15]
port 575 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 wbs_dat_o[16]
port 576 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 wbs_dat_o[17]
port 577 nsew signal output
rlabel metal2 s 37830 0 37886 800 6 wbs_dat_o[18]
port 578 nsew signal output
rlabel metal2 s 39578 0 39634 800 6 wbs_dat_o[19]
port 579 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_o[1]
port 580 nsew signal output
rlabel metal2 s 41326 0 41382 800 6 wbs_dat_o[20]
port 581 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 wbs_dat_o[21]
port 582 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 wbs_dat_o[22]
port 583 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 wbs_dat_o[23]
port 584 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 wbs_dat_o[24]
port 585 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 wbs_dat_o[25]
port 586 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 wbs_dat_o[26]
port 587 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 wbs_dat_o[27]
port 588 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 wbs_dat_o[28]
port 589 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 wbs_dat_o[29]
port 590 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 wbs_dat_o[2]
port 591 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 wbs_dat_o[30]
port 592 nsew signal output
rlabel metal2 s 60094 0 60150 800 6 wbs_dat_o[31]
port 593 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_o[3]
port 594 nsew signal output
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_o[4]
port 595 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_o[5]
port 596 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_o[6]
port 597 nsew signal output
rlabel metal2 s 19062 0 19118 800 6 wbs_dat_o[7]
port 598 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_o[8]
port 599 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 wbs_dat_o[9]
port 600 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 wbs_sel_i[0]
port 601 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wbs_sel_i[1]
port 602 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_sel_i[2]
port 603 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_sel_i[3]
port 604 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_stb_i
port 605 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_we_i
port 606 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 279315 281459
string LEFview TRUE
string GDS_FILE /project/openlane/accelerator_top/runs/accelerator_top/results/magic/accelerator_top.gds
string GDS_END 154754060
string GDS_START 1379770
<< end >>

