magic
tech sky130A
magscale 1 2
timestamp 1636734240
<< obsli1 >>
rect 1104 1377 271308 272017
<< obsm1 >>
rect 14 1300 272214 272048
<< metal2 >>
rect 1122 273827 1178 274627
rect 3422 273827 3478 274627
rect 5814 273827 5870 274627
rect 8206 273827 8262 274627
rect 10598 273827 10654 274627
rect 12990 273827 13046 274627
rect 15382 273827 15438 274627
rect 17774 273827 17830 274627
rect 20166 273827 20222 274627
rect 22558 273827 22614 274627
rect 24950 273827 25006 274627
rect 27342 273827 27398 274627
rect 29734 273827 29790 274627
rect 32126 273827 32182 274627
rect 34518 273827 34574 274627
rect 36910 273827 36966 274627
rect 39302 273827 39358 274627
rect 41694 273827 41750 274627
rect 44086 273827 44142 274627
rect 46478 273827 46534 274627
rect 48870 273827 48926 274627
rect 51262 273827 51318 274627
rect 53654 273827 53710 274627
rect 56046 273827 56102 274627
rect 58438 273827 58494 274627
rect 60830 273827 60886 274627
rect 63222 273827 63278 274627
rect 65614 273827 65670 274627
rect 68006 273827 68062 274627
rect 70398 273827 70454 274627
rect 72790 273827 72846 274627
rect 75182 273827 75238 274627
rect 77574 273827 77630 274627
rect 79966 273827 80022 274627
rect 82358 273827 82414 274627
rect 84750 273827 84806 274627
rect 87142 273827 87198 274627
rect 89534 273827 89590 274627
rect 91926 273827 91982 274627
rect 94318 273827 94374 274627
rect 96710 273827 96766 274627
rect 99102 273827 99158 274627
rect 101494 273827 101550 274627
rect 103886 273827 103942 274627
rect 106278 273827 106334 274627
rect 108670 273827 108726 274627
rect 111062 273827 111118 274627
rect 113454 273827 113510 274627
rect 115846 273827 115902 274627
rect 118238 273827 118294 274627
rect 120630 273827 120686 274627
rect 123022 273827 123078 274627
rect 125414 273827 125470 274627
rect 127806 273827 127862 274627
rect 130198 273827 130254 274627
rect 132590 273827 132646 274627
rect 134982 273827 135038 274627
rect 137374 273827 137430 274627
rect 139674 273827 139730 274627
rect 142066 273827 142122 274627
rect 144458 273827 144514 274627
rect 146850 273827 146906 274627
rect 149242 273827 149298 274627
rect 151634 273827 151690 274627
rect 154026 273827 154082 274627
rect 156418 273827 156474 274627
rect 158810 273827 158866 274627
rect 161202 273827 161258 274627
rect 163594 273827 163650 274627
rect 165986 273827 166042 274627
rect 168378 273827 168434 274627
rect 170770 273827 170826 274627
rect 173162 273827 173218 274627
rect 175554 273827 175610 274627
rect 177946 273827 178002 274627
rect 180338 273827 180394 274627
rect 182730 273827 182786 274627
rect 185122 273827 185178 274627
rect 187514 273827 187570 274627
rect 189906 273827 189962 274627
rect 192298 273827 192354 274627
rect 194690 273827 194746 274627
rect 197082 273827 197138 274627
rect 199474 273827 199530 274627
rect 201866 273827 201922 274627
rect 204258 273827 204314 274627
rect 206650 273827 206706 274627
rect 209042 273827 209098 274627
rect 211434 273827 211490 274627
rect 213826 273827 213882 274627
rect 216218 273827 216274 274627
rect 218610 273827 218666 274627
rect 221002 273827 221058 274627
rect 223394 273827 223450 274627
rect 225786 273827 225842 274627
rect 228178 273827 228234 274627
rect 230570 273827 230626 274627
rect 232962 273827 233018 274627
rect 235354 273827 235410 274627
rect 237746 273827 237802 274627
rect 240138 273827 240194 274627
rect 242530 273827 242586 274627
rect 244922 273827 244978 274627
rect 247314 273827 247370 274627
rect 249706 273827 249762 274627
rect 252098 273827 252154 274627
rect 254490 273827 254546 274627
rect 256882 273827 256938 274627
rect 259274 273827 259330 274627
rect 261666 273827 261722 274627
rect 264058 273827 264114 274627
rect 266450 273827 266506 274627
rect 268842 273827 268898 274627
rect 271234 273827 271290 274627
rect 294 0 350 800
rect 846 0 902 800
rect 1398 0 1454 800
rect 1950 0 2006 800
rect 2502 0 2558 800
rect 3054 0 3110 800
rect 3606 0 3662 800
rect 4158 0 4214 800
rect 4710 0 4766 800
rect 5262 0 5318 800
rect 5814 0 5870 800
rect 6366 0 6422 800
rect 6918 0 6974 800
rect 7470 0 7526 800
rect 8022 0 8078 800
rect 8574 0 8630 800
rect 9126 0 9182 800
rect 9678 0 9734 800
rect 10230 0 10286 800
rect 10782 0 10838 800
rect 11334 0 11390 800
rect 11886 0 11942 800
rect 12438 0 12494 800
rect 13082 0 13138 800
rect 13634 0 13690 800
rect 14186 0 14242 800
rect 14738 0 14794 800
rect 15290 0 15346 800
rect 15842 0 15898 800
rect 16394 0 16450 800
rect 16946 0 17002 800
rect 17498 0 17554 800
rect 18050 0 18106 800
rect 18602 0 18658 800
rect 19154 0 19210 800
rect 19706 0 19762 800
rect 20258 0 20314 800
rect 20810 0 20866 800
rect 21362 0 21418 800
rect 21914 0 21970 800
rect 22466 0 22522 800
rect 23018 0 23074 800
rect 23570 0 23626 800
rect 24122 0 24178 800
rect 24674 0 24730 800
rect 25318 0 25374 800
rect 25870 0 25926 800
rect 26422 0 26478 800
rect 26974 0 27030 800
rect 27526 0 27582 800
rect 28078 0 28134 800
rect 28630 0 28686 800
rect 29182 0 29238 800
rect 29734 0 29790 800
rect 30286 0 30342 800
rect 30838 0 30894 800
rect 31390 0 31446 800
rect 31942 0 31998 800
rect 32494 0 32550 800
rect 33046 0 33102 800
rect 33598 0 33654 800
rect 34150 0 34206 800
rect 34702 0 34758 800
rect 35254 0 35310 800
rect 35806 0 35862 800
rect 36358 0 36414 800
rect 36910 0 36966 800
rect 37554 0 37610 800
rect 38106 0 38162 800
rect 38658 0 38714 800
rect 39210 0 39266 800
rect 39762 0 39818 800
rect 40314 0 40370 800
rect 40866 0 40922 800
rect 41418 0 41474 800
rect 41970 0 42026 800
rect 42522 0 42578 800
rect 43074 0 43130 800
rect 43626 0 43682 800
rect 44178 0 44234 800
rect 44730 0 44786 800
rect 45282 0 45338 800
rect 45834 0 45890 800
rect 46386 0 46442 800
rect 46938 0 46994 800
rect 47490 0 47546 800
rect 48042 0 48098 800
rect 48594 0 48650 800
rect 49146 0 49202 800
rect 49698 0 49754 800
rect 50342 0 50398 800
rect 50894 0 50950 800
rect 51446 0 51502 800
rect 51998 0 52054 800
rect 52550 0 52606 800
rect 53102 0 53158 800
rect 53654 0 53710 800
rect 54206 0 54262 800
rect 54758 0 54814 800
rect 55310 0 55366 800
rect 55862 0 55918 800
rect 56414 0 56470 800
rect 56966 0 57022 800
rect 57518 0 57574 800
rect 58070 0 58126 800
rect 58622 0 58678 800
rect 59174 0 59230 800
rect 59726 0 59782 800
rect 60278 0 60334 800
rect 60830 0 60886 800
rect 61382 0 61438 800
rect 61934 0 61990 800
rect 62578 0 62634 800
rect 63130 0 63186 800
rect 63682 0 63738 800
rect 64234 0 64290 800
rect 64786 0 64842 800
rect 65338 0 65394 800
rect 65890 0 65946 800
rect 66442 0 66498 800
rect 66994 0 67050 800
rect 67546 0 67602 800
rect 68098 0 68154 800
rect 68650 0 68706 800
rect 69202 0 69258 800
rect 69754 0 69810 800
rect 70306 0 70362 800
rect 70858 0 70914 800
rect 71410 0 71466 800
rect 71962 0 72018 800
rect 72514 0 72570 800
rect 73066 0 73122 800
rect 73618 0 73674 800
rect 74170 0 74226 800
rect 74814 0 74870 800
rect 75366 0 75422 800
rect 75918 0 75974 800
rect 76470 0 76526 800
rect 77022 0 77078 800
rect 77574 0 77630 800
rect 78126 0 78182 800
rect 78678 0 78734 800
rect 79230 0 79286 800
rect 79782 0 79838 800
rect 80334 0 80390 800
rect 80886 0 80942 800
rect 81438 0 81494 800
rect 81990 0 82046 800
rect 82542 0 82598 800
rect 83094 0 83150 800
rect 83646 0 83702 800
rect 84198 0 84254 800
rect 84750 0 84806 800
rect 85302 0 85358 800
rect 85854 0 85910 800
rect 86406 0 86462 800
rect 87050 0 87106 800
rect 87602 0 87658 800
rect 88154 0 88210 800
rect 88706 0 88762 800
rect 89258 0 89314 800
rect 89810 0 89866 800
rect 90362 0 90418 800
rect 90914 0 90970 800
rect 91466 0 91522 800
rect 92018 0 92074 800
rect 92570 0 92626 800
rect 93122 0 93178 800
rect 93674 0 93730 800
rect 94226 0 94282 800
rect 94778 0 94834 800
rect 95330 0 95386 800
rect 95882 0 95938 800
rect 96434 0 96490 800
rect 96986 0 97042 800
rect 97538 0 97594 800
rect 98090 0 98146 800
rect 98642 0 98698 800
rect 99194 0 99250 800
rect 99838 0 99894 800
rect 100390 0 100446 800
rect 100942 0 100998 800
rect 101494 0 101550 800
rect 102046 0 102102 800
rect 102598 0 102654 800
rect 103150 0 103206 800
rect 103702 0 103758 800
rect 104254 0 104310 800
rect 104806 0 104862 800
rect 105358 0 105414 800
rect 105910 0 105966 800
rect 106462 0 106518 800
rect 107014 0 107070 800
rect 107566 0 107622 800
rect 108118 0 108174 800
rect 108670 0 108726 800
rect 109222 0 109278 800
rect 109774 0 109830 800
rect 110326 0 110382 800
rect 110878 0 110934 800
rect 111430 0 111486 800
rect 112074 0 112130 800
rect 112626 0 112682 800
rect 113178 0 113234 800
rect 113730 0 113786 800
rect 114282 0 114338 800
rect 114834 0 114890 800
rect 115386 0 115442 800
rect 115938 0 115994 800
rect 116490 0 116546 800
rect 117042 0 117098 800
rect 117594 0 117650 800
rect 118146 0 118202 800
rect 118698 0 118754 800
rect 119250 0 119306 800
rect 119802 0 119858 800
rect 120354 0 120410 800
rect 120906 0 120962 800
rect 121458 0 121514 800
rect 122010 0 122066 800
rect 122562 0 122618 800
rect 123114 0 123170 800
rect 123666 0 123722 800
rect 124310 0 124366 800
rect 124862 0 124918 800
rect 125414 0 125470 800
rect 125966 0 126022 800
rect 126518 0 126574 800
rect 127070 0 127126 800
rect 127622 0 127678 800
rect 128174 0 128230 800
rect 128726 0 128782 800
rect 129278 0 129334 800
rect 129830 0 129886 800
rect 130382 0 130438 800
rect 130934 0 130990 800
rect 131486 0 131542 800
rect 132038 0 132094 800
rect 132590 0 132646 800
rect 133142 0 133198 800
rect 133694 0 133750 800
rect 134246 0 134302 800
rect 134798 0 134854 800
rect 135350 0 135406 800
rect 135902 0 135958 800
rect 136546 0 136602 800
rect 137098 0 137154 800
rect 137650 0 137706 800
rect 138202 0 138258 800
rect 138754 0 138810 800
rect 139306 0 139362 800
rect 139858 0 139914 800
rect 140410 0 140466 800
rect 140962 0 141018 800
rect 141514 0 141570 800
rect 142066 0 142122 800
rect 142618 0 142674 800
rect 143170 0 143226 800
rect 143722 0 143778 800
rect 144274 0 144330 800
rect 144826 0 144882 800
rect 145378 0 145434 800
rect 145930 0 145986 800
rect 146482 0 146538 800
rect 147034 0 147090 800
rect 147586 0 147642 800
rect 148138 0 148194 800
rect 148690 0 148746 800
rect 149334 0 149390 800
rect 149886 0 149942 800
rect 150438 0 150494 800
rect 150990 0 151046 800
rect 151542 0 151598 800
rect 152094 0 152150 800
rect 152646 0 152702 800
rect 153198 0 153254 800
rect 153750 0 153806 800
rect 154302 0 154358 800
rect 154854 0 154910 800
rect 155406 0 155462 800
rect 155958 0 156014 800
rect 156510 0 156566 800
rect 157062 0 157118 800
rect 157614 0 157670 800
rect 158166 0 158222 800
rect 158718 0 158774 800
rect 159270 0 159326 800
rect 159822 0 159878 800
rect 160374 0 160430 800
rect 160926 0 160982 800
rect 161570 0 161626 800
rect 162122 0 162178 800
rect 162674 0 162730 800
rect 163226 0 163282 800
rect 163778 0 163834 800
rect 164330 0 164386 800
rect 164882 0 164938 800
rect 165434 0 165490 800
rect 165986 0 166042 800
rect 166538 0 166594 800
rect 167090 0 167146 800
rect 167642 0 167698 800
rect 168194 0 168250 800
rect 168746 0 168802 800
rect 169298 0 169354 800
rect 169850 0 169906 800
rect 170402 0 170458 800
rect 170954 0 171010 800
rect 171506 0 171562 800
rect 172058 0 172114 800
rect 172610 0 172666 800
rect 173162 0 173218 800
rect 173806 0 173862 800
rect 174358 0 174414 800
rect 174910 0 174966 800
rect 175462 0 175518 800
rect 176014 0 176070 800
rect 176566 0 176622 800
rect 177118 0 177174 800
rect 177670 0 177726 800
rect 178222 0 178278 800
rect 178774 0 178830 800
rect 179326 0 179382 800
rect 179878 0 179934 800
rect 180430 0 180486 800
rect 180982 0 181038 800
rect 181534 0 181590 800
rect 182086 0 182142 800
rect 182638 0 182694 800
rect 183190 0 183246 800
rect 183742 0 183798 800
rect 184294 0 184350 800
rect 184846 0 184902 800
rect 185398 0 185454 800
rect 185950 0 186006 800
rect 186594 0 186650 800
rect 187146 0 187202 800
rect 187698 0 187754 800
rect 188250 0 188306 800
rect 188802 0 188858 800
rect 189354 0 189410 800
rect 189906 0 189962 800
rect 190458 0 190514 800
rect 191010 0 191066 800
rect 191562 0 191618 800
rect 192114 0 192170 800
rect 192666 0 192722 800
rect 193218 0 193274 800
rect 193770 0 193826 800
rect 194322 0 194378 800
rect 194874 0 194930 800
rect 195426 0 195482 800
rect 195978 0 196034 800
rect 196530 0 196586 800
rect 197082 0 197138 800
rect 197634 0 197690 800
rect 198186 0 198242 800
rect 198830 0 198886 800
rect 199382 0 199438 800
rect 199934 0 199990 800
rect 200486 0 200542 800
rect 201038 0 201094 800
rect 201590 0 201646 800
rect 202142 0 202198 800
rect 202694 0 202750 800
rect 203246 0 203302 800
rect 203798 0 203854 800
rect 204350 0 204406 800
rect 204902 0 204958 800
rect 205454 0 205510 800
rect 206006 0 206062 800
rect 206558 0 206614 800
rect 207110 0 207166 800
rect 207662 0 207718 800
rect 208214 0 208270 800
rect 208766 0 208822 800
rect 209318 0 209374 800
rect 209870 0 209926 800
rect 210422 0 210478 800
rect 211066 0 211122 800
rect 211618 0 211674 800
rect 212170 0 212226 800
rect 212722 0 212778 800
rect 213274 0 213330 800
rect 213826 0 213882 800
rect 214378 0 214434 800
rect 214930 0 214986 800
rect 215482 0 215538 800
rect 216034 0 216090 800
rect 216586 0 216642 800
rect 217138 0 217194 800
rect 217690 0 217746 800
rect 218242 0 218298 800
rect 218794 0 218850 800
rect 219346 0 219402 800
rect 219898 0 219954 800
rect 220450 0 220506 800
rect 221002 0 221058 800
rect 221554 0 221610 800
rect 222106 0 222162 800
rect 222658 0 222714 800
rect 223302 0 223358 800
rect 223854 0 223910 800
rect 224406 0 224462 800
rect 224958 0 225014 800
rect 225510 0 225566 800
rect 226062 0 226118 800
rect 226614 0 226670 800
rect 227166 0 227222 800
rect 227718 0 227774 800
rect 228270 0 228326 800
rect 228822 0 228878 800
rect 229374 0 229430 800
rect 229926 0 229982 800
rect 230478 0 230534 800
rect 231030 0 231086 800
rect 231582 0 231638 800
rect 232134 0 232190 800
rect 232686 0 232742 800
rect 233238 0 233294 800
rect 233790 0 233846 800
rect 234342 0 234398 800
rect 234894 0 234950 800
rect 235446 0 235502 800
rect 236090 0 236146 800
rect 236642 0 236698 800
rect 237194 0 237250 800
rect 237746 0 237802 800
rect 238298 0 238354 800
rect 238850 0 238906 800
rect 239402 0 239458 800
rect 239954 0 240010 800
rect 240506 0 240562 800
rect 241058 0 241114 800
rect 241610 0 241666 800
rect 242162 0 242218 800
rect 242714 0 242770 800
rect 243266 0 243322 800
rect 243818 0 243874 800
rect 244370 0 244426 800
rect 244922 0 244978 800
rect 245474 0 245530 800
rect 246026 0 246082 800
rect 246578 0 246634 800
rect 247130 0 247186 800
rect 247682 0 247738 800
rect 248326 0 248382 800
rect 248878 0 248934 800
rect 249430 0 249486 800
rect 249982 0 250038 800
rect 250534 0 250590 800
rect 251086 0 251142 800
rect 251638 0 251694 800
rect 252190 0 252246 800
rect 252742 0 252798 800
rect 253294 0 253350 800
rect 253846 0 253902 800
rect 254398 0 254454 800
rect 254950 0 255006 800
rect 255502 0 255558 800
rect 256054 0 256110 800
rect 256606 0 256662 800
rect 257158 0 257214 800
rect 257710 0 257766 800
rect 258262 0 258318 800
rect 258814 0 258870 800
rect 259366 0 259422 800
rect 259918 0 259974 800
rect 260562 0 260618 800
rect 261114 0 261170 800
rect 261666 0 261722 800
rect 262218 0 262274 800
rect 262770 0 262826 800
rect 263322 0 263378 800
rect 263874 0 263930 800
rect 264426 0 264482 800
rect 264978 0 265034 800
rect 265530 0 265586 800
rect 266082 0 266138 800
rect 266634 0 266690 800
rect 267186 0 267242 800
rect 267738 0 267794 800
rect 268290 0 268346 800
rect 268842 0 268898 800
rect 269394 0 269450 800
rect 269946 0 270002 800
rect 270498 0 270554 800
rect 271050 0 271106 800
rect 271602 0 271658 800
rect 272154 0 272210 800
<< obsm2 >>
rect 20 273771 1066 273827
rect 1234 273771 3366 273827
rect 3534 273771 5758 273827
rect 5926 273771 8150 273827
rect 8318 273771 10542 273827
rect 10710 273771 12934 273827
rect 13102 273771 15326 273827
rect 15494 273771 17718 273827
rect 17886 273771 20110 273827
rect 20278 273771 22502 273827
rect 22670 273771 24894 273827
rect 25062 273771 27286 273827
rect 27454 273771 29678 273827
rect 29846 273771 32070 273827
rect 32238 273771 34462 273827
rect 34630 273771 36854 273827
rect 37022 273771 39246 273827
rect 39414 273771 41638 273827
rect 41806 273771 44030 273827
rect 44198 273771 46422 273827
rect 46590 273771 48814 273827
rect 48982 273771 51206 273827
rect 51374 273771 53598 273827
rect 53766 273771 55990 273827
rect 56158 273771 58382 273827
rect 58550 273771 60774 273827
rect 60942 273771 63166 273827
rect 63334 273771 65558 273827
rect 65726 273771 67950 273827
rect 68118 273771 70342 273827
rect 70510 273771 72734 273827
rect 72902 273771 75126 273827
rect 75294 273771 77518 273827
rect 77686 273771 79910 273827
rect 80078 273771 82302 273827
rect 82470 273771 84694 273827
rect 84862 273771 87086 273827
rect 87254 273771 89478 273827
rect 89646 273771 91870 273827
rect 92038 273771 94262 273827
rect 94430 273771 96654 273827
rect 96822 273771 99046 273827
rect 99214 273771 101438 273827
rect 101606 273771 103830 273827
rect 103998 273771 106222 273827
rect 106390 273771 108614 273827
rect 108782 273771 111006 273827
rect 111174 273771 113398 273827
rect 113566 273771 115790 273827
rect 115958 273771 118182 273827
rect 118350 273771 120574 273827
rect 120742 273771 122966 273827
rect 123134 273771 125358 273827
rect 125526 273771 127750 273827
rect 127918 273771 130142 273827
rect 130310 273771 132534 273827
rect 132702 273771 134926 273827
rect 135094 273771 137318 273827
rect 137486 273771 139618 273827
rect 139786 273771 142010 273827
rect 142178 273771 144402 273827
rect 144570 273771 146794 273827
rect 146962 273771 149186 273827
rect 149354 273771 151578 273827
rect 151746 273771 153970 273827
rect 154138 273771 156362 273827
rect 156530 273771 158754 273827
rect 158922 273771 161146 273827
rect 161314 273771 163538 273827
rect 163706 273771 165930 273827
rect 166098 273771 168322 273827
rect 168490 273771 170714 273827
rect 170882 273771 173106 273827
rect 173274 273771 175498 273827
rect 175666 273771 177890 273827
rect 178058 273771 180282 273827
rect 180450 273771 182674 273827
rect 182842 273771 185066 273827
rect 185234 273771 187458 273827
rect 187626 273771 189850 273827
rect 190018 273771 192242 273827
rect 192410 273771 194634 273827
rect 194802 273771 197026 273827
rect 197194 273771 199418 273827
rect 199586 273771 201810 273827
rect 201978 273771 204202 273827
rect 204370 273771 206594 273827
rect 206762 273771 208986 273827
rect 209154 273771 211378 273827
rect 211546 273771 213770 273827
rect 213938 273771 216162 273827
rect 216330 273771 218554 273827
rect 218722 273771 220946 273827
rect 221114 273771 223338 273827
rect 223506 273771 225730 273827
rect 225898 273771 228122 273827
rect 228290 273771 230514 273827
rect 230682 273771 232906 273827
rect 233074 273771 235298 273827
rect 235466 273771 237690 273827
rect 237858 273771 240082 273827
rect 240250 273771 242474 273827
rect 242642 273771 244866 273827
rect 245034 273771 247258 273827
rect 247426 273771 249650 273827
rect 249818 273771 252042 273827
rect 252210 273771 254434 273827
rect 254602 273771 256826 273827
rect 256994 273771 259218 273827
rect 259386 273771 261610 273827
rect 261778 273771 264002 273827
rect 264170 273771 266394 273827
rect 266562 273771 268786 273827
rect 268954 273771 271178 273827
rect 271346 273771 272208 273827
rect 20 856 272208 273771
rect 20 734 238 856
rect 406 734 790 856
rect 958 734 1342 856
rect 1510 734 1894 856
rect 2062 734 2446 856
rect 2614 734 2998 856
rect 3166 734 3550 856
rect 3718 734 4102 856
rect 4270 734 4654 856
rect 4822 734 5206 856
rect 5374 734 5758 856
rect 5926 734 6310 856
rect 6478 734 6862 856
rect 7030 734 7414 856
rect 7582 734 7966 856
rect 8134 734 8518 856
rect 8686 734 9070 856
rect 9238 734 9622 856
rect 9790 734 10174 856
rect 10342 734 10726 856
rect 10894 734 11278 856
rect 11446 734 11830 856
rect 11998 734 12382 856
rect 12550 734 13026 856
rect 13194 734 13578 856
rect 13746 734 14130 856
rect 14298 734 14682 856
rect 14850 734 15234 856
rect 15402 734 15786 856
rect 15954 734 16338 856
rect 16506 734 16890 856
rect 17058 734 17442 856
rect 17610 734 17994 856
rect 18162 734 18546 856
rect 18714 734 19098 856
rect 19266 734 19650 856
rect 19818 734 20202 856
rect 20370 734 20754 856
rect 20922 734 21306 856
rect 21474 734 21858 856
rect 22026 734 22410 856
rect 22578 734 22962 856
rect 23130 734 23514 856
rect 23682 734 24066 856
rect 24234 734 24618 856
rect 24786 734 25262 856
rect 25430 734 25814 856
rect 25982 734 26366 856
rect 26534 734 26918 856
rect 27086 734 27470 856
rect 27638 734 28022 856
rect 28190 734 28574 856
rect 28742 734 29126 856
rect 29294 734 29678 856
rect 29846 734 30230 856
rect 30398 734 30782 856
rect 30950 734 31334 856
rect 31502 734 31886 856
rect 32054 734 32438 856
rect 32606 734 32990 856
rect 33158 734 33542 856
rect 33710 734 34094 856
rect 34262 734 34646 856
rect 34814 734 35198 856
rect 35366 734 35750 856
rect 35918 734 36302 856
rect 36470 734 36854 856
rect 37022 734 37498 856
rect 37666 734 38050 856
rect 38218 734 38602 856
rect 38770 734 39154 856
rect 39322 734 39706 856
rect 39874 734 40258 856
rect 40426 734 40810 856
rect 40978 734 41362 856
rect 41530 734 41914 856
rect 42082 734 42466 856
rect 42634 734 43018 856
rect 43186 734 43570 856
rect 43738 734 44122 856
rect 44290 734 44674 856
rect 44842 734 45226 856
rect 45394 734 45778 856
rect 45946 734 46330 856
rect 46498 734 46882 856
rect 47050 734 47434 856
rect 47602 734 47986 856
rect 48154 734 48538 856
rect 48706 734 49090 856
rect 49258 734 49642 856
rect 49810 734 50286 856
rect 50454 734 50838 856
rect 51006 734 51390 856
rect 51558 734 51942 856
rect 52110 734 52494 856
rect 52662 734 53046 856
rect 53214 734 53598 856
rect 53766 734 54150 856
rect 54318 734 54702 856
rect 54870 734 55254 856
rect 55422 734 55806 856
rect 55974 734 56358 856
rect 56526 734 56910 856
rect 57078 734 57462 856
rect 57630 734 58014 856
rect 58182 734 58566 856
rect 58734 734 59118 856
rect 59286 734 59670 856
rect 59838 734 60222 856
rect 60390 734 60774 856
rect 60942 734 61326 856
rect 61494 734 61878 856
rect 62046 734 62522 856
rect 62690 734 63074 856
rect 63242 734 63626 856
rect 63794 734 64178 856
rect 64346 734 64730 856
rect 64898 734 65282 856
rect 65450 734 65834 856
rect 66002 734 66386 856
rect 66554 734 66938 856
rect 67106 734 67490 856
rect 67658 734 68042 856
rect 68210 734 68594 856
rect 68762 734 69146 856
rect 69314 734 69698 856
rect 69866 734 70250 856
rect 70418 734 70802 856
rect 70970 734 71354 856
rect 71522 734 71906 856
rect 72074 734 72458 856
rect 72626 734 73010 856
rect 73178 734 73562 856
rect 73730 734 74114 856
rect 74282 734 74758 856
rect 74926 734 75310 856
rect 75478 734 75862 856
rect 76030 734 76414 856
rect 76582 734 76966 856
rect 77134 734 77518 856
rect 77686 734 78070 856
rect 78238 734 78622 856
rect 78790 734 79174 856
rect 79342 734 79726 856
rect 79894 734 80278 856
rect 80446 734 80830 856
rect 80998 734 81382 856
rect 81550 734 81934 856
rect 82102 734 82486 856
rect 82654 734 83038 856
rect 83206 734 83590 856
rect 83758 734 84142 856
rect 84310 734 84694 856
rect 84862 734 85246 856
rect 85414 734 85798 856
rect 85966 734 86350 856
rect 86518 734 86994 856
rect 87162 734 87546 856
rect 87714 734 88098 856
rect 88266 734 88650 856
rect 88818 734 89202 856
rect 89370 734 89754 856
rect 89922 734 90306 856
rect 90474 734 90858 856
rect 91026 734 91410 856
rect 91578 734 91962 856
rect 92130 734 92514 856
rect 92682 734 93066 856
rect 93234 734 93618 856
rect 93786 734 94170 856
rect 94338 734 94722 856
rect 94890 734 95274 856
rect 95442 734 95826 856
rect 95994 734 96378 856
rect 96546 734 96930 856
rect 97098 734 97482 856
rect 97650 734 98034 856
rect 98202 734 98586 856
rect 98754 734 99138 856
rect 99306 734 99782 856
rect 99950 734 100334 856
rect 100502 734 100886 856
rect 101054 734 101438 856
rect 101606 734 101990 856
rect 102158 734 102542 856
rect 102710 734 103094 856
rect 103262 734 103646 856
rect 103814 734 104198 856
rect 104366 734 104750 856
rect 104918 734 105302 856
rect 105470 734 105854 856
rect 106022 734 106406 856
rect 106574 734 106958 856
rect 107126 734 107510 856
rect 107678 734 108062 856
rect 108230 734 108614 856
rect 108782 734 109166 856
rect 109334 734 109718 856
rect 109886 734 110270 856
rect 110438 734 110822 856
rect 110990 734 111374 856
rect 111542 734 112018 856
rect 112186 734 112570 856
rect 112738 734 113122 856
rect 113290 734 113674 856
rect 113842 734 114226 856
rect 114394 734 114778 856
rect 114946 734 115330 856
rect 115498 734 115882 856
rect 116050 734 116434 856
rect 116602 734 116986 856
rect 117154 734 117538 856
rect 117706 734 118090 856
rect 118258 734 118642 856
rect 118810 734 119194 856
rect 119362 734 119746 856
rect 119914 734 120298 856
rect 120466 734 120850 856
rect 121018 734 121402 856
rect 121570 734 121954 856
rect 122122 734 122506 856
rect 122674 734 123058 856
rect 123226 734 123610 856
rect 123778 734 124254 856
rect 124422 734 124806 856
rect 124974 734 125358 856
rect 125526 734 125910 856
rect 126078 734 126462 856
rect 126630 734 127014 856
rect 127182 734 127566 856
rect 127734 734 128118 856
rect 128286 734 128670 856
rect 128838 734 129222 856
rect 129390 734 129774 856
rect 129942 734 130326 856
rect 130494 734 130878 856
rect 131046 734 131430 856
rect 131598 734 131982 856
rect 132150 734 132534 856
rect 132702 734 133086 856
rect 133254 734 133638 856
rect 133806 734 134190 856
rect 134358 734 134742 856
rect 134910 734 135294 856
rect 135462 734 135846 856
rect 136014 734 136490 856
rect 136658 734 137042 856
rect 137210 734 137594 856
rect 137762 734 138146 856
rect 138314 734 138698 856
rect 138866 734 139250 856
rect 139418 734 139802 856
rect 139970 734 140354 856
rect 140522 734 140906 856
rect 141074 734 141458 856
rect 141626 734 142010 856
rect 142178 734 142562 856
rect 142730 734 143114 856
rect 143282 734 143666 856
rect 143834 734 144218 856
rect 144386 734 144770 856
rect 144938 734 145322 856
rect 145490 734 145874 856
rect 146042 734 146426 856
rect 146594 734 146978 856
rect 147146 734 147530 856
rect 147698 734 148082 856
rect 148250 734 148634 856
rect 148802 734 149278 856
rect 149446 734 149830 856
rect 149998 734 150382 856
rect 150550 734 150934 856
rect 151102 734 151486 856
rect 151654 734 152038 856
rect 152206 734 152590 856
rect 152758 734 153142 856
rect 153310 734 153694 856
rect 153862 734 154246 856
rect 154414 734 154798 856
rect 154966 734 155350 856
rect 155518 734 155902 856
rect 156070 734 156454 856
rect 156622 734 157006 856
rect 157174 734 157558 856
rect 157726 734 158110 856
rect 158278 734 158662 856
rect 158830 734 159214 856
rect 159382 734 159766 856
rect 159934 734 160318 856
rect 160486 734 160870 856
rect 161038 734 161514 856
rect 161682 734 162066 856
rect 162234 734 162618 856
rect 162786 734 163170 856
rect 163338 734 163722 856
rect 163890 734 164274 856
rect 164442 734 164826 856
rect 164994 734 165378 856
rect 165546 734 165930 856
rect 166098 734 166482 856
rect 166650 734 167034 856
rect 167202 734 167586 856
rect 167754 734 168138 856
rect 168306 734 168690 856
rect 168858 734 169242 856
rect 169410 734 169794 856
rect 169962 734 170346 856
rect 170514 734 170898 856
rect 171066 734 171450 856
rect 171618 734 172002 856
rect 172170 734 172554 856
rect 172722 734 173106 856
rect 173274 734 173750 856
rect 173918 734 174302 856
rect 174470 734 174854 856
rect 175022 734 175406 856
rect 175574 734 175958 856
rect 176126 734 176510 856
rect 176678 734 177062 856
rect 177230 734 177614 856
rect 177782 734 178166 856
rect 178334 734 178718 856
rect 178886 734 179270 856
rect 179438 734 179822 856
rect 179990 734 180374 856
rect 180542 734 180926 856
rect 181094 734 181478 856
rect 181646 734 182030 856
rect 182198 734 182582 856
rect 182750 734 183134 856
rect 183302 734 183686 856
rect 183854 734 184238 856
rect 184406 734 184790 856
rect 184958 734 185342 856
rect 185510 734 185894 856
rect 186062 734 186538 856
rect 186706 734 187090 856
rect 187258 734 187642 856
rect 187810 734 188194 856
rect 188362 734 188746 856
rect 188914 734 189298 856
rect 189466 734 189850 856
rect 190018 734 190402 856
rect 190570 734 190954 856
rect 191122 734 191506 856
rect 191674 734 192058 856
rect 192226 734 192610 856
rect 192778 734 193162 856
rect 193330 734 193714 856
rect 193882 734 194266 856
rect 194434 734 194818 856
rect 194986 734 195370 856
rect 195538 734 195922 856
rect 196090 734 196474 856
rect 196642 734 197026 856
rect 197194 734 197578 856
rect 197746 734 198130 856
rect 198298 734 198774 856
rect 198942 734 199326 856
rect 199494 734 199878 856
rect 200046 734 200430 856
rect 200598 734 200982 856
rect 201150 734 201534 856
rect 201702 734 202086 856
rect 202254 734 202638 856
rect 202806 734 203190 856
rect 203358 734 203742 856
rect 203910 734 204294 856
rect 204462 734 204846 856
rect 205014 734 205398 856
rect 205566 734 205950 856
rect 206118 734 206502 856
rect 206670 734 207054 856
rect 207222 734 207606 856
rect 207774 734 208158 856
rect 208326 734 208710 856
rect 208878 734 209262 856
rect 209430 734 209814 856
rect 209982 734 210366 856
rect 210534 734 211010 856
rect 211178 734 211562 856
rect 211730 734 212114 856
rect 212282 734 212666 856
rect 212834 734 213218 856
rect 213386 734 213770 856
rect 213938 734 214322 856
rect 214490 734 214874 856
rect 215042 734 215426 856
rect 215594 734 215978 856
rect 216146 734 216530 856
rect 216698 734 217082 856
rect 217250 734 217634 856
rect 217802 734 218186 856
rect 218354 734 218738 856
rect 218906 734 219290 856
rect 219458 734 219842 856
rect 220010 734 220394 856
rect 220562 734 220946 856
rect 221114 734 221498 856
rect 221666 734 222050 856
rect 222218 734 222602 856
rect 222770 734 223246 856
rect 223414 734 223798 856
rect 223966 734 224350 856
rect 224518 734 224902 856
rect 225070 734 225454 856
rect 225622 734 226006 856
rect 226174 734 226558 856
rect 226726 734 227110 856
rect 227278 734 227662 856
rect 227830 734 228214 856
rect 228382 734 228766 856
rect 228934 734 229318 856
rect 229486 734 229870 856
rect 230038 734 230422 856
rect 230590 734 230974 856
rect 231142 734 231526 856
rect 231694 734 232078 856
rect 232246 734 232630 856
rect 232798 734 233182 856
rect 233350 734 233734 856
rect 233902 734 234286 856
rect 234454 734 234838 856
rect 235006 734 235390 856
rect 235558 734 236034 856
rect 236202 734 236586 856
rect 236754 734 237138 856
rect 237306 734 237690 856
rect 237858 734 238242 856
rect 238410 734 238794 856
rect 238962 734 239346 856
rect 239514 734 239898 856
rect 240066 734 240450 856
rect 240618 734 241002 856
rect 241170 734 241554 856
rect 241722 734 242106 856
rect 242274 734 242658 856
rect 242826 734 243210 856
rect 243378 734 243762 856
rect 243930 734 244314 856
rect 244482 734 244866 856
rect 245034 734 245418 856
rect 245586 734 245970 856
rect 246138 734 246522 856
rect 246690 734 247074 856
rect 247242 734 247626 856
rect 247794 734 248270 856
rect 248438 734 248822 856
rect 248990 734 249374 856
rect 249542 734 249926 856
rect 250094 734 250478 856
rect 250646 734 251030 856
rect 251198 734 251582 856
rect 251750 734 252134 856
rect 252302 734 252686 856
rect 252854 734 253238 856
rect 253406 734 253790 856
rect 253958 734 254342 856
rect 254510 734 254894 856
rect 255062 734 255446 856
rect 255614 734 255998 856
rect 256166 734 256550 856
rect 256718 734 257102 856
rect 257270 734 257654 856
rect 257822 734 258206 856
rect 258374 734 258758 856
rect 258926 734 259310 856
rect 259478 734 259862 856
rect 260030 734 260506 856
rect 260674 734 261058 856
rect 261226 734 261610 856
rect 261778 734 262162 856
rect 262330 734 262714 856
rect 262882 734 263266 856
rect 263434 734 263818 856
rect 263986 734 264370 856
rect 264538 734 264922 856
rect 265090 734 265474 856
rect 265642 734 266026 856
rect 266194 734 266578 856
rect 266746 734 267130 856
rect 267298 734 267682 856
rect 267850 734 268234 856
rect 268402 734 268786 856
rect 268954 734 269338 856
rect 269506 734 269890 856
rect 270058 734 270442 856
rect 270610 734 270994 856
rect 271162 734 271546 856
rect 271714 734 272098 856
<< obsm3 >>
rect 3049 2143 265648 272033
<< metal4 >>
rect 4208 2128 4528 272048
rect 19568 2128 19888 272048
rect 34928 2128 35248 272048
rect 50288 2128 50608 272048
rect 65648 2128 65968 272048
rect 81008 2128 81328 272048
rect 96368 2128 96688 272048
rect 111728 2128 112048 272048
rect 127088 2128 127408 272048
rect 142448 2128 142768 272048
rect 157808 2128 158128 272048
rect 173168 2128 173488 272048
rect 188528 2128 188848 272048
rect 203888 2128 204208 272048
rect 219248 2128 219568 272048
rect 234608 2128 234928 272048
rect 249968 2128 250288 272048
rect 265328 2128 265648 272048
<< obsm4 >>
rect 3923 2619 4128 260133
rect 4608 2619 19488 260133
rect 19968 2619 34848 260133
rect 35328 2619 50208 260133
rect 50688 2619 65568 260133
rect 66048 2619 80928 260133
rect 81408 2619 96288 260133
rect 96768 2619 111648 260133
rect 112128 2619 127008 260133
rect 127488 2619 142368 260133
rect 142848 2619 157728 260133
rect 158208 2619 173088 260133
rect 173568 2619 188448 260133
rect 188928 2619 203808 260133
rect 204288 2619 219168 260133
rect 219648 2619 221109 260133
<< labels >>
rlabel metal2 s 1122 273827 1178 274627 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 72790 273827 72846 274627 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 79966 273827 80022 274627 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 87142 273827 87198 274627 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 94318 273827 94374 274627 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 101494 273827 101550 274627 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 108670 273827 108726 274627 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 115846 273827 115902 274627 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 123022 273827 123078 274627 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 130198 273827 130254 274627 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 137374 273827 137430 274627 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 8206 273827 8262 274627 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 144458 273827 144514 274627 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 151634 273827 151690 274627 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 158810 273827 158866 274627 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 165986 273827 166042 274627 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 173162 273827 173218 274627 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 180338 273827 180394 274627 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 187514 273827 187570 274627 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 194690 273827 194746 274627 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 201866 273827 201922 274627 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 209042 273827 209098 274627 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 15382 273827 15438 274627 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 216218 273827 216274 274627 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 223394 273827 223450 274627 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 230570 273827 230626 274627 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 237746 273827 237802 274627 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 244922 273827 244978 274627 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 252098 273827 252154 274627 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 259274 273827 259330 274627 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 266450 273827 266506 274627 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 22558 273827 22614 274627 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 29734 273827 29790 274627 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 36910 273827 36966 274627 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 44086 273827 44142 274627 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 51262 273827 51318 274627 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 58438 273827 58494 274627 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 65614 273827 65670 274627 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3422 273827 3478 274627 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 75182 273827 75238 274627 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 82358 273827 82414 274627 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 89534 273827 89590 274627 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 96710 273827 96766 274627 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 103886 273827 103942 274627 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 111062 273827 111118 274627 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 118238 273827 118294 274627 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 125414 273827 125470 274627 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 132590 273827 132646 274627 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 139674 273827 139730 274627 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 10598 273827 10654 274627 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 146850 273827 146906 274627 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 154026 273827 154082 274627 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 161202 273827 161258 274627 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 168378 273827 168434 274627 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 175554 273827 175610 274627 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 182730 273827 182786 274627 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 189906 273827 189962 274627 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 197082 273827 197138 274627 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 204258 273827 204314 274627 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 211434 273827 211490 274627 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 17774 273827 17830 274627 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 218610 273827 218666 274627 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 225786 273827 225842 274627 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 232962 273827 233018 274627 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 240138 273827 240194 274627 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 247314 273827 247370 274627 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 254490 273827 254546 274627 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 261666 273827 261722 274627 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 268842 273827 268898 274627 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 24950 273827 25006 274627 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 32126 273827 32182 274627 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 39302 273827 39358 274627 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 46478 273827 46534 274627 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 53654 273827 53710 274627 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 60830 273827 60886 274627 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 68006 273827 68062 274627 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 5814 273827 5870 274627 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 77574 273827 77630 274627 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 84750 273827 84806 274627 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 91926 273827 91982 274627 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 99102 273827 99158 274627 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 106278 273827 106334 274627 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 113454 273827 113510 274627 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 120630 273827 120686 274627 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 127806 273827 127862 274627 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 134982 273827 135038 274627 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 142066 273827 142122 274627 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 12990 273827 13046 274627 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 149242 273827 149298 274627 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 156418 273827 156474 274627 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 163594 273827 163650 274627 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 170770 273827 170826 274627 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 177946 273827 178002 274627 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 185122 273827 185178 274627 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 192298 273827 192354 274627 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 199474 273827 199530 274627 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 206650 273827 206706 274627 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 213826 273827 213882 274627 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 20166 273827 20222 274627 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 221002 273827 221058 274627 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 228178 273827 228234 274627 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 235354 273827 235410 274627 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 242530 273827 242586 274627 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 249706 273827 249762 274627 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 256882 273827 256938 274627 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 264058 273827 264114 274627 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 271234 273827 271290 274627 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 27342 273827 27398 274627 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 34518 273827 34574 274627 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 41694 273827 41750 274627 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 48870 273827 48926 274627 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 56046 273827 56102 274627 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 63222 273827 63278 274627 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 70398 273827 70454 274627 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 59174 0 59230 800 6 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 226062 0 226118 800 6 la_data_in[100]
port 116 nsew signal input
rlabel metal2 s 227718 0 227774 800 6 la_data_in[101]
port 117 nsew signal input
rlabel metal2 s 229374 0 229430 800 6 la_data_in[102]
port 118 nsew signal input
rlabel metal2 s 231030 0 231086 800 6 la_data_in[103]
port 119 nsew signal input
rlabel metal2 s 232686 0 232742 800 6 la_data_in[104]
port 120 nsew signal input
rlabel metal2 s 234342 0 234398 800 6 la_data_in[105]
port 121 nsew signal input
rlabel metal2 s 236090 0 236146 800 6 la_data_in[106]
port 122 nsew signal input
rlabel metal2 s 237746 0 237802 800 6 la_data_in[107]
port 123 nsew signal input
rlabel metal2 s 239402 0 239458 800 6 la_data_in[108]
port 124 nsew signal input
rlabel metal2 s 241058 0 241114 800 6 la_data_in[109]
port 125 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_data_in[10]
port 126 nsew signal input
rlabel metal2 s 242714 0 242770 800 6 la_data_in[110]
port 127 nsew signal input
rlabel metal2 s 244370 0 244426 800 6 la_data_in[111]
port 128 nsew signal input
rlabel metal2 s 246026 0 246082 800 6 la_data_in[112]
port 129 nsew signal input
rlabel metal2 s 247682 0 247738 800 6 la_data_in[113]
port 130 nsew signal input
rlabel metal2 s 249430 0 249486 800 6 la_data_in[114]
port 131 nsew signal input
rlabel metal2 s 251086 0 251142 800 6 la_data_in[115]
port 132 nsew signal input
rlabel metal2 s 252742 0 252798 800 6 la_data_in[116]
port 133 nsew signal input
rlabel metal2 s 254398 0 254454 800 6 la_data_in[117]
port 134 nsew signal input
rlabel metal2 s 256054 0 256110 800 6 la_data_in[118]
port 135 nsew signal input
rlabel metal2 s 257710 0 257766 800 6 la_data_in[119]
port 136 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_data_in[11]
port 137 nsew signal input
rlabel metal2 s 259366 0 259422 800 6 la_data_in[120]
port 138 nsew signal input
rlabel metal2 s 261114 0 261170 800 6 la_data_in[121]
port 139 nsew signal input
rlabel metal2 s 262770 0 262826 800 6 la_data_in[122]
port 140 nsew signal input
rlabel metal2 s 264426 0 264482 800 6 la_data_in[123]
port 141 nsew signal input
rlabel metal2 s 266082 0 266138 800 6 la_data_in[124]
port 142 nsew signal input
rlabel metal2 s 267738 0 267794 800 6 la_data_in[125]
port 143 nsew signal input
rlabel metal2 s 269394 0 269450 800 6 la_data_in[126]
port 144 nsew signal input
rlabel metal2 s 271050 0 271106 800 6 la_data_in[127]
port 145 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_data_in[12]
port 146 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 la_data_in[13]
port 147 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_data_in[14]
port 148 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_data_in[15]
port 149 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_data_in[16]
port 150 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 la_data_in[17]
port 151 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 la_data_in[18]
port 152 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_data_in[19]
port 153 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 la_data_in[1]
port 154 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_data_in[20]
port 155 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_data_in[21]
port 156 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 la_data_in[22]
port 157 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 la_data_in[23]
port 158 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_data_in[24]
port 159 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 la_data_in[25]
port 160 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 la_data_in[26]
port 161 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 la_data_in[27]
port 162 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 la_data_in[28]
port 163 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_data_in[29]
port 164 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 la_data_in[2]
port 165 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 la_data_in[30]
port 166 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 la_data_in[31]
port 167 nsew signal input
rlabel metal2 s 112626 0 112682 800 6 la_data_in[32]
port 168 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 la_data_in[33]
port 169 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 la_data_in[34]
port 170 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 la_data_in[35]
port 171 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 la_data_in[36]
port 172 nsew signal input
rlabel metal2 s 120906 0 120962 800 6 la_data_in[37]
port 173 nsew signal input
rlabel metal2 s 122562 0 122618 800 6 la_data_in[38]
port 174 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 la_data_in[39]
port 175 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 la_data_in[3]
port 176 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 la_data_in[40]
port 177 nsew signal input
rlabel metal2 s 127622 0 127678 800 6 la_data_in[41]
port 178 nsew signal input
rlabel metal2 s 129278 0 129334 800 6 la_data_in[42]
port 179 nsew signal input
rlabel metal2 s 130934 0 130990 800 6 la_data_in[43]
port 180 nsew signal input
rlabel metal2 s 132590 0 132646 800 6 la_data_in[44]
port 181 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 la_data_in[45]
port 182 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 la_data_in[46]
port 183 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 la_data_in[47]
port 184 nsew signal input
rlabel metal2 s 139306 0 139362 800 6 la_data_in[48]
port 185 nsew signal input
rlabel metal2 s 140962 0 141018 800 6 la_data_in[49]
port 186 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 la_data_in[4]
port 187 nsew signal input
rlabel metal2 s 142618 0 142674 800 6 la_data_in[50]
port 188 nsew signal input
rlabel metal2 s 144274 0 144330 800 6 la_data_in[51]
port 189 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 la_data_in[52]
port 190 nsew signal input
rlabel metal2 s 147586 0 147642 800 6 la_data_in[53]
port 191 nsew signal input
rlabel metal2 s 149334 0 149390 800 6 la_data_in[54]
port 192 nsew signal input
rlabel metal2 s 150990 0 151046 800 6 la_data_in[55]
port 193 nsew signal input
rlabel metal2 s 152646 0 152702 800 6 la_data_in[56]
port 194 nsew signal input
rlabel metal2 s 154302 0 154358 800 6 la_data_in[57]
port 195 nsew signal input
rlabel metal2 s 155958 0 156014 800 6 la_data_in[58]
port 196 nsew signal input
rlabel metal2 s 157614 0 157670 800 6 la_data_in[59]
port 197 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_data_in[5]
port 198 nsew signal input
rlabel metal2 s 159270 0 159326 800 6 la_data_in[60]
port 199 nsew signal input
rlabel metal2 s 160926 0 160982 800 6 la_data_in[61]
port 200 nsew signal input
rlabel metal2 s 162674 0 162730 800 6 la_data_in[62]
port 201 nsew signal input
rlabel metal2 s 164330 0 164386 800 6 la_data_in[63]
port 202 nsew signal input
rlabel metal2 s 165986 0 166042 800 6 la_data_in[64]
port 203 nsew signal input
rlabel metal2 s 167642 0 167698 800 6 la_data_in[65]
port 204 nsew signal input
rlabel metal2 s 169298 0 169354 800 6 la_data_in[66]
port 205 nsew signal input
rlabel metal2 s 170954 0 171010 800 6 la_data_in[67]
port 206 nsew signal input
rlabel metal2 s 172610 0 172666 800 6 la_data_in[68]
port 207 nsew signal input
rlabel metal2 s 174358 0 174414 800 6 la_data_in[69]
port 208 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_data_in[6]
port 209 nsew signal input
rlabel metal2 s 176014 0 176070 800 6 la_data_in[70]
port 210 nsew signal input
rlabel metal2 s 177670 0 177726 800 6 la_data_in[71]
port 211 nsew signal input
rlabel metal2 s 179326 0 179382 800 6 la_data_in[72]
port 212 nsew signal input
rlabel metal2 s 180982 0 181038 800 6 la_data_in[73]
port 213 nsew signal input
rlabel metal2 s 182638 0 182694 800 6 la_data_in[74]
port 214 nsew signal input
rlabel metal2 s 184294 0 184350 800 6 la_data_in[75]
port 215 nsew signal input
rlabel metal2 s 185950 0 186006 800 6 la_data_in[76]
port 216 nsew signal input
rlabel metal2 s 187698 0 187754 800 6 la_data_in[77]
port 217 nsew signal input
rlabel metal2 s 189354 0 189410 800 6 la_data_in[78]
port 218 nsew signal input
rlabel metal2 s 191010 0 191066 800 6 la_data_in[79]
port 219 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 la_data_in[7]
port 220 nsew signal input
rlabel metal2 s 192666 0 192722 800 6 la_data_in[80]
port 221 nsew signal input
rlabel metal2 s 194322 0 194378 800 6 la_data_in[81]
port 222 nsew signal input
rlabel metal2 s 195978 0 196034 800 6 la_data_in[82]
port 223 nsew signal input
rlabel metal2 s 197634 0 197690 800 6 la_data_in[83]
port 224 nsew signal input
rlabel metal2 s 199382 0 199438 800 6 la_data_in[84]
port 225 nsew signal input
rlabel metal2 s 201038 0 201094 800 6 la_data_in[85]
port 226 nsew signal input
rlabel metal2 s 202694 0 202750 800 6 la_data_in[86]
port 227 nsew signal input
rlabel metal2 s 204350 0 204406 800 6 la_data_in[87]
port 228 nsew signal input
rlabel metal2 s 206006 0 206062 800 6 la_data_in[88]
port 229 nsew signal input
rlabel metal2 s 207662 0 207718 800 6 la_data_in[89]
port 230 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 la_data_in[8]
port 231 nsew signal input
rlabel metal2 s 209318 0 209374 800 6 la_data_in[90]
port 232 nsew signal input
rlabel metal2 s 211066 0 211122 800 6 la_data_in[91]
port 233 nsew signal input
rlabel metal2 s 212722 0 212778 800 6 la_data_in[92]
port 234 nsew signal input
rlabel metal2 s 214378 0 214434 800 6 la_data_in[93]
port 235 nsew signal input
rlabel metal2 s 216034 0 216090 800 6 la_data_in[94]
port 236 nsew signal input
rlabel metal2 s 217690 0 217746 800 6 la_data_in[95]
port 237 nsew signal input
rlabel metal2 s 219346 0 219402 800 6 la_data_in[96]
port 238 nsew signal input
rlabel metal2 s 221002 0 221058 800 6 la_data_in[97]
port 239 nsew signal input
rlabel metal2 s 222658 0 222714 800 6 la_data_in[98]
port 240 nsew signal input
rlabel metal2 s 224406 0 224462 800 6 la_data_in[99]
port 241 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 la_data_in[9]
port 242 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 la_data_out[0]
port 243 nsew signal output
rlabel metal2 s 226614 0 226670 800 6 la_data_out[100]
port 244 nsew signal output
rlabel metal2 s 228270 0 228326 800 6 la_data_out[101]
port 245 nsew signal output
rlabel metal2 s 229926 0 229982 800 6 la_data_out[102]
port 246 nsew signal output
rlabel metal2 s 231582 0 231638 800 6 la_data_out[103]
port 247 nsew signal output
rlabel metal2 s 233238 0 233294 800 6 la_data_out[104]
port 248 nsew signal output
rlabel metal2 s 234894 0 234950 800 6 la_data_out[105]
port 249 nsew signal output
rlabel metal2 s 236642 0 236698 800 6 la_data_out[106]
port 250 nsew signal output
rlabel metal2 s 238298 0 238354 800 6 la_data_out[107]
port 251 nsew signal output
rlabel metal2 s 239954 0 240010 800 6 la_data_out[108]
port 252 nsew signal output
rlabel metal2 s 241610 0 241666 800 6 la_data_out[109]
port 253 nsew signal output
rlabel metal2 s 76470 0 76526 800 6 la_data_out[10]
port 254 nsew signal output
rlabel metal2 s 243266 0 243322 800 6 la_data_out[110]
port 255 nsew signal output
rlabel metal2 s 244922 0 244978 800 6 la_data_out[111]
port 256 nsew signal output
rlabel metal2 s 246578 0 246634 800 6 la_data_out[112]
port 257 nsew signal output
rlabel metal2 s 248326 0 248382 800 6 la_data_out[113]
port 258 nsew signal output
rlabel metal2 s 249982 0 250038 800 6 la_data_out[114]
port 259 nsew signal output
rlabel metal2 s 251638 0 251694 800 6 la_data_out[115]
port 260 nsew signal output
rlabel metal2 s 253294 0 253350 800 6 la_data_out[116]
port 261 nsew signal output
rlabel metal2 s 254950 0 255006 800 6 la_data_out[117]
port 262 nsew signal output
rlabel metal2 s 256606 0 256662 800 6 la_data_out[118]
port 263 nsew signal output
rlabel metal2 s 258262 0 258318 800 6 la_data_out[119]
port 264 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 la_data_out[11]
port 265 nsew signal output
rlabel metal2 s 259918 0 259974 800 6 la_data_out[120]
port 266 nsew signal output
rlabel metal2 s 261666 0 261722 800 6 la_data_out[121]
port 267 nsew signal output
rlabel metal2 s 263322 0 263378 800 6 la_data_out[122]
port 268 nsew signal output
rlabel metal2 s 264978 0 265034 800 6 la_data_out[123]
port 269 nsew signal output
rlabel metal2 s 266634 0 266690 800 6 la_data_out[124]
port 270 nsew signal output
rlabel metal2 s 268290 0 268346 800 6 la_data_out[125]
port 271 nsew signal output
rlabel metal2 s 269946 0 270002 800 6 la_data_out[126]
port 272 nsew signal output
rlabel metal2 s 271602 0 271658 800 6 la_data_out[127]
port 273 nsew signal output
rlabel metal2 s 79782 0 79838 800 6 la_data_out[12]
port 274 nsew signal output
rlabel metal2 s 81438 0 81494 800 6 la_data_out[13]
port 275 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 la_data_out[14]
port 276 nsew signal output
rlabel metal2 s 84750 0 84806 800 6 la_data_out[15]
port 277 nsew signal output
rlabel metal2 s 86406 0 86462 800 6 la_data_out[16]
port 278 nsew signal output
rlabel metal2 s 88154 0 88210 800 6 la_data_out[17]
port 279 nsew signal output
rlabel metal2 s 89810 0 89866 800 6 la_data_out[18]
port 280 nsew signal output
rlabel metal2 s 91466 0 91522 800 6 la_data_out[19]
port 281 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 la_data_out[1]
port 282 nsew signal output
rlabel metal2 s 93122 0 93178 800 6 la_data_out[20]
port 283 nsew signal output
rlabel metal2 s 94778 0 94834 800 6 la_data_out[21]
port 284 nsew signal output
rlabel metal2 s 96434 0 96490 800 6 la_data_out[22]
port 285 nsew signal output
rlabel metal2 s 98090 0 98146 800 6 la_data_out[23]
port 286 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 la_data_out[24]
port 287 nsew signal output
rlabel metal2 s 101494 0 101550 800 6 la_data_out[25]
port 288 nsew signal output
rlabel metal2 s 103150 0 103206 800 6 la_data_out[26]
port 289 nsew signal output
rlabel metal2 s 104806 0 104862 800 6 la_data_out[27]
port 290 nsew signal output
rlabel metal2 s 106462 0 106518 800 6 la_data_out[28]
port 291 nsew signal output
rlabel metal2 s 108118 0 108174 800 6 la_data_out[29]
port 292 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 la_data_out[2]
port 293 nsew signal output
rlabel metal2 s 109774 0 109830 800 6 la_data_out[30]
port 294 nsew signal output
rlabel metal2 s 111430 0 111486 800 6 la_data_out[31]
port 295 nsew signal output
rlabel metal2 s 113178 0 113234 800 6 la_data_out[32]
port 296 nsew signal output
rlabel metal2 s 114834 0 114890 800 6 la_data_out[33]
port 297 nsew signal output
rlabel metal2 s 116490 0 116546 800 6 la_data_out[34]
port 298 nsew signal output
rlabel metal2 s 118146 0 118202 800 6 la_data_out[35]
port 299 nsew signal output
rlabel metal2 s 119802 0 119858 800 6 la_data_out[36]
port 300 nsew signal output
rlabel metal2 s 121458 0 121514 800 6 la_data_out[37]
port 301 nsew signal output
rlabel metal2 s 123114 0 123170 800 6 la_data_out[38]
port 302 nsew signal output
rlabel metal2 s 124862 0 124918 800 6 la_data_out[39]
port 303 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 la_data_out[3]
port 304 nsew signal output
rlabel metal2 s 126518 0 126574 800 6 la_data_out[40]
port 305 nsew signal output
rlabel metal2 s 128174 0 128230 800 6 la_data_out[41]
port 306 nsew signal output
rlabel metal2 s 129830 0 129886 800 6 la_data_out[42]
port 307 nsew signal output
rlabel metal2 s 131486 0 131542 800 6 la_data_out[43]
port 308 nsew signal output
rlabel metal2 s 133142 0 133198 800 6 la_data_out[44]
port 309 nsew signal output
rlabel metal2 s 134798 0 134854 800 6 la_data_out[45]
port 310 nsew signal output
rlabel metal2 s 136546 0 136602 800 6 la_data_out[46]
port 311 nsew signal output
rlabel metal2 s 138202 0 138258 800 6 la_data_out[47]
port 312 nsew signal output
rlabel metal2 s 139858 0 139914 800 6 la_data_out[48]
port 313 nsew signal output
rlabel metal2 s 141514 0 141570 800 6 la_data_out[49]
port 314 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 la_data_out[4]
port 315 nsew signal output
rlabel metal2 s 143170 0 143226 800 6 la_data_out[50]
port 316 nsew signal output
rlabel metal2 s 144826 0 144882 800 6 la_data_out[51]
port 317 nsew signal output
rlabel metal2 s 146482 0 146538 800 6 la_data_out[52]
port 318 nsew signal output
rlabel metal2 s 148138 0 148194 800 6 la_data_out[53]
port 319 nsew signal output
rlabel metal2 s 149886 0 149942 800 6 la_data_out[54]
port 320 nsew signal output
rlabel metal2 s 151542 0 151598 800 6 la_data_out[55]
port 321 nsew signal output
rlabel metal2 s 153198 0 153254 800 6 la_data_out[56]
port 322 nsew signal output
rlabel metal2 s 154854 0 154910 800 6 la_data_out[57]
port 323 nsew signal output
rlabel metal2 s 156510 0 156566 800 6 la_data_out[58]
port 324 nsew signal output
rlabel metal2 s 158166 0 158222 800 6 la_data_out[59]
port 325 nsew signal output
rlabel metal2 s 68098 0 68154 800 6 la_data_out[5]
port 326 nsew signal output
rlabel metal2 s 159822 0 159878 800 6 la_data_out[60]
port 327 nsew signal output
rlabel metal2 s 161570 0 161626 800 6 la_data_out[61]
port 328 nsew signal output
rlabel metal2 s 163226 0 163282 800 6 la_data_out[62]
port 329 nsew signal output
rlabel metal2 s 164882 0 164938 800 6 la_data_out[63]
port 330 nsew signal output
rlabel metal2 s 166538 0 166594 800 6 la_data_out[64]
port 331 nsew signal output
rlabel metal2 s 168194 0 168250 800 6 la_data_out[65]
port 332 nsew signal output
rlabel metal2 s 169850 0 169906 800 6 la_data_out[66]
port 333 nsew signal output
rlabel metal2 s 171506 0 171562 800 6 la_data_out[67]
port 334 nsew signal output
rlabel metal2 s 173162 0 173218 800 6 la_data_out[68]
port 335 nsew signal output
rlabel metal2 s 174910 0 174966 800 6 la_data_out[69]
port 336 nsew signal output
rlabel metal2 s 69754 0 69810 800 6 la_data_out[6]
port 337 nsew signal output
rlabel metal2 s 176566 0 176622 800 6 la_data_out[70]
port 338 nsew signal output
rlabel metal2 s 178222 0 178278 800 6 la_data_out[71]
port 339 nsew signal output
rlabel metal2 s 179878 0 179934 800 6 la_data_out[72]
port 340 nsew signal output
rlabel metal2 s 181534 0 181590 800 6 la_data_out[73]
port 341 nsew signal output
rlabel metal2 s 183190 0 183246 800 6 la_data_out[74]
port 342 nsew signal output
rlabel metal2 s 184846 0 184902 800 6 la_data_out[75]
port 343 nsew signal output
rlabel metal2 s 186594 0 186650 800 6 la_data_out[76]
port 344 nsew signal output
rlabel metal2 s 188250 0 188306 800 6 la_data_out[77]
port 345 nsew signal output
rlabel metal2 s 189906 0 189962 800 6 la_data_out[78]
port 346 nsew signal output
rlabel metal2 s 191562 0 191618 800 6 la_data_out[79]
port 347 nsew signal output
rlabel metal2 s 71410 0 71466 800 6 la_data_out[7]
port 348 nsew signal output
rlabel metal2 s 193218 0 193274 800 6 la_data_out[80]
port 349 nsew signal output
rlabel metal2 s 194874 0 194930 800 6 la_data_out[81]
port 350 nsew signal output
rlabel metal2 s 196530 0 196586 800 6 la_data_out[82]
port 351 nsew signal output
rlabel metal2 s 198186 0 198242 800 6 la_data_out[83]
port 352 nsew signal output
rlabel metal2 s 199934 0 199990 800 6 la_data_out[84]
port 353 nsew signal output
rlabel metal2 s 201590 0 201646 800 6 la_data_out[85]
port 354 nsew signal output
rlabel metal2 s 203246 0 203302 800 6 la_data_out[86]
port 355 nsew signal output
rlabel metal2 s 204902 0 204958 800 6 la_data_out[87]
port 356 nsew signal output
rlabel metal2 s 206558 0 206614 800 6 la_data_out[88]
port 357 nsew signal output
rlabel metal2 s 208214 0 208270 800 6 la_data_out[89]
port 358 nsew signal output
rlabel metal2 s 73066 0 73122 800 6 la_data_out[8]
port 359 nsew signal output
rlabel metal2 s 209870 0 209926 800 6 la_data_out[90]
port 360 nsew signal output
rlabel metal2 s 211618 0 211674 800 6 la_data_out[91]
port 361 nsew signal output
rlabel metal2 s 213274 0 213330 800 6 la_data_out[92]
port 362 nsew signal output
rlabel metal2 s 214930 0 214986 800 6 la_data_out[93]
port 363 nsew signal output
rlabel metal2 s 216586 0 216642 800 6 la_data_out[94]
port 364 nsew signal output
rlabel metal2 s 218242 0 218298 800 6 la_data_out[95]
port 365 nsew signal output
rlabel metal2 s 219898 0 219954 800 6 la_data_out[96]
port 366 nsew signal output
rlabel metal2 s 221554 0 221610 800 6 la_data_out[97]
port 367 nsew signal output
rlabel metal2 s 223302 0 223358 800 6 la_data_out[98]
port 368 nsew signal output
rlabel metal2 s 224958 0 225014 800 6 la_data_out[99]
port 369 nsew signal output
rlabel metal2 s 74814 0 74870 800 6 la_data_out[9]
port 370 nsew signal output
rlabel metal2 s 60278 0 60334 800 6 la_oen[0]
port 371 nsew signal input
rlabel metal2 s 227166 0 227222 800 6 la_oen[100]
port 372 nsew signal input
rlabel metal2 s 228822 0 228878 800 6 la_oen[101]
port 373 nsew signal input
rlabel metal2 s 230478 0 230534 800 6 la_oen[102]
port 374 nsew signal input
rlabel metal2 s 232134 0 232190 800 6 la_oen[103]
port 375 nsew signal input
rlabel metal2 s 233790 0 233846 800 6 la_oen[104]
port 376 nsew signal input
rlabel metal2 s 235446 0 235502 800 6 la_oen[105]
port 377 nsew signal input
rlabel metal2 s 237194 0 237250 800 6 la_oen[106]
port 378 nsew signal input
rlabel metal2 s 238850 0 238906 800 6 la_oen[107]
port 379 nsew signal input
rlabel metal2 s 240506 0 240562 800 6 la_oen[108]
port 380 nsew signal input
rlabel metal2 s 242162 0 242218 800 6 la_oen[109]
port 381 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 la_oen[10]
port 382 nsew signal input
rlabel metal2 s 243818 0 243874 800 6 la_oen[110]
port 383 nsew signal input
rlabel metal2 s 245474 0 245530 800 6 la_oen[111]
port 384 nsew signal input
rlabel metal2 s 247130 0 247186 800 6 la_oen[112]
port 385 nsew signal input
rlabel metal2 s 248878 0 248934 800 6 la_oen[113]
port 386 nsew signal input
rlabel metal2 s 250534 0 250590 800 6 la_oen[114]
port 387 nsew signal input
rlabel metal2 s 252190 0 252246 800 6 la_oen[115]
port 388 nsew signal input
rlabel metal2 s 253846 0 253902 800 6 la_oen[116]
port 389 nsew signal input
rlabel metal2 s 255502 0 255558 800 6 la_oen[117]
port 390 nsew signal input
rlabel metal2 s 257158 0 257214 800 6 la_oen[118]
port 391 nsew signal input
rlabel metal2 s 258814 0 258870 800 6 la_oen[119]
port 392 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 la_oen[11]
port 393 nsew signal input
rlabel metal2 s 260562 0 260618 800 6 la_oen[120]
port 394 nsew signal input
rlabel metal2 s 262218 0 262274 800 6 la_oen[121]
port 395 nsew signal input
rlabel metal2 s 263874 0 263930 800 6 la_oen[122]
port 396 nsew signal input
rlabel metal2 s 265530 0 265586 800 6 la_oen[123]
port 397 nsew signal input
rlabel metal2 s 267186 0 267242 800 6 la_oen[124]
port 398 nsew signal input
rlabel metal2 s 268842 0 268898 800 6 la_oen[125]
port 399 nsew signal input
rlabel metal2 s 270498 0 270554 800 6 la_oen[126]
port 400 nsew signal input
rlabel metal2 s 272154 0 272210 800 6 la_oen[127]
port 401 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_oen[12]
port 402 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_oen[13]
port 403 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_oen[14]
port 404 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_oen[15]
port 405 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_oen[16]
port 406 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_oen[17]
port 407 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 la_oen[18]
port 408 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_oen[19]
port 409 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 la_oen[1]
port 410 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_oen[20]
port 411 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 la_oen[21]
port 412 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_oen[22]
port 413 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_oen[23]
port 414 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_oen[24]
port 415 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 la_oen[25]
port 416 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_oen[26]
port 417 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 la_oen[27]
port 418 nsew signal input
rlabel metal2 s 107014 0 107070 800 6 la_oen[28]
port 419 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 la_oen[29]
port 420 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 la_oen[2]
port 421 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 la_oen[30]
port 422 nsew signal input
rlabel metal2 s 112074 0 112130 800 6 la_oen[31]
port 423 nsew signal input
rlabel metal2 s 113730 0 113786 800 6 la_oen[32]
port 424 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 la_oen[33]
port 425 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 la_oen[34]
port 426 nsew signal input
rlabel metal2 s 118698 0 118754 800 6 la_oen[35]
port 427 nsew signal input
rlabel metal2 s 120354 0 120410 800 6 la_oen[36]
port 428 nsew signal input
rlabel metal2 s 122010 0 122066 800 6 la_oen[37]
port 429 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 la_oen[38]
port 430 nsew signal input
rlabel metal2 s 125414 0 125470 800 6 la_oen[39]
port 431 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_oen[3]
port 432 nsew signal input
rlabel metal2 s 127070 0 127126 800 6 la_oen[40]
port 433 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 la_oen[41]
port 434 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 la_oen[42]
port 435 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 la_oen[43]
port 436 nsew signal input
rlabel metal2 s 133694 0 133750 800 6 la_oen[44]
port 437 nsew signal input
rlabel metal2 s 135350 0 135406 800 6 la_oen[45]
port 438 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 la_oen[46]
port 439 nsew signal input
rlabel metal2 s 138754 0 138810 800 6 la_oen[47]
port 440 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_oen[48]
port 441 nsew signal input
rlabel metal2 s 142066 0 142122 800 6 la_oen[49]
port 442 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 la_oen[4]
port 443 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 la_oen[50]
port 444 nsew signal input
rlabel metal2 s 145378 0 145434 800 6 la_oen[51]
port 445 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 la_oen[52]
port 446 nsew signal input
rlabel metal2 s 148690 0 148746 800 6 la_oen[53]
port 447 nsew signal input
rlabel metal2 s 150438 0 150494 800 6 la_oen[54]
port 448 nsew signal input
rlabel metal2 s 152094 0 152150 800 6 la_oen[55]
port 449 nsew signal input
rlabel metal2 s 153750 0 153806 800 6 la_oen[56]
port 450 nsew signal input
rlabel metal2 s 155406 0 155462 800 6 la_oen[57]
port 451 nsew signal input
rlabel metal2 s 157062 0 157118 800 6 la_oen[58]
port 452 nsew signal input
rlabel metal2 s 158718 0 158774 800 6 la_oen[59]
port 453 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 la_oen[5]
port 454 nsew signal input
rlabel metal2 s 160374 0 160430 800 6 la_oen[60]
port 455 nsew signal input
rlabel metal2 s 162122 0 162178 800 6 la_oen[61]
port 456 nsew signal input
rlabel metal2 s 163778 0 163834 800 6 la_oen[62]
port 457 nsew signal input
rlabel metal2 s 165434 0 165490 800 6 la_oen[63]
port 458 nsew signal input
rlabel metal2 s 167090 0 167146 800 6 la_oen[64]
port 459 nsew signal input
rlabel metal2 s 168746 0 168802 800 6 la_oen[65]
port 460 nsew signal input
rlabel metal2 s 170402 0 170458 800 6 la_oen[66]
port 461 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 la_oen[67]
port 462 nsew signal input
rlabel metal2 s 173806 0 173862 800 6 la_oen[68]
port 463 nsew signal input
rlabel metal2 s 175462 0 175518 800 6 la_oen[69]
port 464 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 la_oen[6]
port 465 nsew signal input
rlabel metal2 s 177118 0 177174 800 6 la_oen[70]
port 466 nsew signal input
rlabel metal2 s 178774 0 178830 800 6 la_oen[71]
port 467 nsew signal input
rlabel metal2 s 180430 0 180486 800 6 la_oen[72]
port 468 nsew signal input
rlabel metal2 s 182086 0 182142 800 6 la_oen[73]
port 469 nsew signal input
rlabel metal2 s 183742 0 183798 800 6 la_oen[74]
port 470 nsew signal input
rlabel metal2 s 185398 0 185454 800 6 la_oen[75]
port 471 nsew signal input
rlabel metal2 s 187146 0 187202 800 6 la_oen[76]
port 472 nsew signal input
rlabel metal2 s 188802 0 188858 800 6 la_oen[77]
port 473 nsew signal input
rlabel metal2 s 190458 0 190514 800 6 la_oen[78]
port 474 nsew signal input
rlabel metal2 s 192114 0 192170 800 6 la_oen[79]
port 475 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 la_oen[7]
port 476 nsew signal input
rlabel metal2 s 193770 0 193826 800 6 la_oen[80]
port 477 nsew signal input
rlabel metal2 s 195426 0 195482 800 6 la_oen[81]
port 478 nsew signal input
rlabel metal2 s 197082 0 197138 800 6 la_oen[82]
port 479 nsew signal input
rlabel metal2 s 198830 0 198886 800 6 la_oen[83]
port 480 nsew signal input
rlabel metal2 s 200486 0 200542 800 6 la_oen[84]
port 481 nsew signal input
rlabel metal2 s 202142 0 202198 800 6 la_oen[85]
port 482 nsew signal input
rlabel metal2 s 203798 0 203854 800 6 la_oen[86]
port 483 nsew signal input
rlabel metal2 s 205454 0 205510 800 6 la_oen[87]
port 484 nsew signal input
rlabel metal2 s 207110 0 207166 800 6 la_oen[88]
port 485 nsew signal input
rlabel metal2 s 208766 0 208822 800 6 la_oen[89]
port 486 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_oen[8]
port 487 nsew signal input
rlabel metal2 s 210422 0 210478 800 6 la_oen[90]
port 488 nsew signal input
rlabel metal2 s 212170 0 212226 800 6 la_oen[91]
port 489 nsew signal input
rlabel metal2 s 213826 0 213882 800 6 la_oen[92]
port 490 nsew signal input
rlabel metal2 s 215482 0 215538 800 6 la_oen[93]
port 491 nsew signal input
rlabel metal2 s 217138 0 217194 800 6 la_oen[94]
port 492 nsew signal input
rlabel metal2 s 218794 0 218850 800 6 la_oen[95]
port 493 nsew signal input
rlabel metal2 s 220450 0 220506 800 6 la_oen[96]
port 494 nsew signal input
rlabel metal2 s 222106 0 222162 800 6 la_oen[97]
port 495 nsew signal input
rlabel metal2 s 223854 0 223910 800 6 la_oen[98]
port 496 nsew signal input
rlabel metal2 s 225510 0 225566 800 6 la_oen[99]
port 497 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_oen[9]
port 498 nsew signal input
rlabel metal4 s 4208 2128 4528 272048 6 vccd1
port 499 nsew power input
rlabel metal4 s 34928 2128 35248 272048 6 vccd1
port 499 nsew power input
rlabel metal4 s 65648 2128 65968 272048 6 vccd1
port 499 nsew power input
rlabel metal4 s 96368 2128 96688 272048 6 vccd1
port 499 nsew power input
rlabel metal4 s 127088 2128 127408 272048 6 vccd1
port 499 nsew power input
rlabel metal4 s 157808 2128 158128 272048 6 vccd1
port 499 nsew power input
rlabel metal4 s 188528 2128 188848 272048 6 vccd1
port 499 nsew power input
rlabel metal4 s 219248 2128 219568 272048 6 vccd1
port 499 nsew power input
rlabel metal4 s 249968 2128 250288 272048 6 vccd1
port 499 nsew power input
rlabel metal4 s 19568 2128 19888 272048 6 vssd1
port 500 nsew ground input
rlabel metal4 s 50288 2128 50608 272048 6 vssd1
port 500 nsew ground input
rlabel metal4 s 81008 2128 81328 272048 6 vssd1
port 500 nsew ground input
rlabel metal4 s 111728 2128 112048 272048 6 vssd1
port 500 nsew ground input
rlabel metal4 s 142448 2128 142768 272048 6 vssd1
port 500 nsew ground input
rlabel metal4 s 173168 2128 173488 272048 6 vssd1
port 500 nsew ground input
rlabel metal4 s 203888 2128 204208 272048 6 vssd1
port 500 nsew ground input
rlabel metal4 s 234608 2128 234928 272048 6 vssd1
port 500 nsew ground input
rlabel metal4 s 265328 2128 265648 272048 6 vssd1
port 500 nsew ground input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 501 nsew signal input
rlabel metal2 s 846 0 902 800 6 wb_rst_i
port 502 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_ack_o
port 503 nsew signal output
rlabel metal2 s 3606 0 3662 800 6 wbs_adr_i[0]
port 504 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_adr_i[10]
port 505 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_adr_i[11]
port 506 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 wbs_adr_i[12]
port 507 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_adr_i[13]
port 508 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wbs_adr_i[14]
port 509 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wbs_adr_i[15]
port 510 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_adr_i[16]
port 511 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 wbs_adr_i[17]
port 512 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 wbs_adr_i[18]
port 513 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 wbs_adr_i[19]
port 514 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_adr_i[1]
port 515 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 wbs_adr_i[20]
port 516 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 wbs_adr_i[21]
port 517 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_adr_i[22]
port 518 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 wbs_adr_i[23]
port 519 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 wbs_adr_i[24]
port 520 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 wbs_adr_i[25]
port 521 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 wbs_adr_i[26]
port 522 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 wbs_adr_i[27]
port 523 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 wbs_adr_i[28]
port 524 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 wbs_adr_i[29]
port 525 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 wbs_adr_i[2]
port 526 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 wbs_adr_i[30]
port 527 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 wbs_adr_i[31]
port 528 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_adr_i[3]
port 529 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_adr_i[4]
port 530 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_adr_i[5]
port 531 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 wbs_adr_i[6]
port 532 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wbs_adr_i[7]
port 533 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_adr_i[8]
port 534 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 wbs_adr_i[9]
port 535 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_cyc_i
port 536 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_dat_i[0]
port 537 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_dat_i[10]
port 538 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_i[11]
port 539 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_i[12]
port 540 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wbs_dat_i[13]
port 541 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_dat_i[14]
port 542 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wbs_dat_i[15]
port 543 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wbs_dat_i[16]
port 544 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 wbs_dat_i[17]
port 545 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wbs_dat_i[18]
port 546 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 wbs_dat_i[19]
port 547 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_dat_i[1]
port 548 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 wbs_dat_i[20]
port 549 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 wbs_dat_i[21]
port 550 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 wbs_dat_i[22]
port 551 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 wbs_dat_i[23]
port 552 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 wbs_dat_i[24]
port 553 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 wbs_dat_i[25]
port 554 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 wbs_dat_i[26]
port 555 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 wbs_dat_i[27]
port 556 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 wbs_dat_i[28]
port 557 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 wbs_dat_i[29]
port 558 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_i[2]
port 559 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 wbs_dat_i[30]
port 560 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 wbs_dat_i[31]
port 561 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_i[3]
port 562 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_i[4]
port 563 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_dat_i[5]
port 564 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_dat_i[6]
port 565 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[7]
port 566 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_i[8]
port 567 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_i[9]
port 568 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_o[0]
port 569 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 wbs_dat_o[10]
port 570 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 wbs_dat_o[11]
port 571 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_o[12]
port 572 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_o[13]
port 573 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_o[14]
port 574 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 wbs_dat_o[15]
port 575 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 wbs_dat_o[16]
port 576 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_o[17]
port 577 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_o[18]
port 578 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_o[19]
port 579 nsew signal output
rlabel metal2 s 6918 0 6974 800 6 wbs_dat_o[1]
port 580 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 wbs_dat_o[20]
port 581 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 wbs_dat_o[21]
port 582 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 wbs_dat_o[22]
port 583 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 wbs_dat_o[23]
port 584 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 wbs_dat_o[24]
port 585 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 wbs_dat_o[25]
port 586 nsew signal output
rlabel metal2 s 50342 0 50398 800 6 wbs_dat_o[26]
port 587 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 wbs_dat_o[27]
port 588 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 wbs_dat_o[28]
port 589 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 wbs_dat_o[29]
port 590 nsew signal output
rlabel metal2 s 9126 0 9182 800 6 wbs_dat_o[2]
port 591 nsew signal output
rlabel metal2 s 56966 0 57022 800 6 wbs_dat_o[30]
port 592 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 wbs_dat_o[31]
port 593 nsew signal output
rlabel metal2 s 11334 0 11390 800 6 wbs_dat_o[3]
port 594 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 wbs_dat_o[4]
port 595 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_o[5]
port 596 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_o[6]
port 597 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_o[7]
port 598 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 wbs_dat_o[8]
port 599 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 wbs_dat_o[9]
port 600 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 wbs_sel_i[0]
port 601 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_sel_i[1]
port 602 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_sel_i[2]
port 603 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_sel_i[3]
port 604 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_stb_i
port 605 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_we_i
port 606 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 272483 274627
string LEFview TRUE
string GDS_FILE /project/openlane/accelerator_top/runs/accelerator_top/results/magic/accelerator_top.gds
string GDS_END 161163876
string GDS_START 1285956
<< end >>

